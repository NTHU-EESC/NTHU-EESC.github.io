************************************************************************
* auCdl Netlist:
* 
* Library Name:  Hw4_3
* Top Cell Name: Differential
* View Name:     schematic
* Netlisted on:  May  7 21:40:17 2015
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: Hw4_3
* Cell Name:    Differential
* View Name:    schematic
************************************************************************

.SUBCKT Differential GND VDD Vin1 Vin2 Vout Vp
*.PININFO GND:I VDD:I Vin1:I Vin2:I Vout:O
MM4 Vout Vx VDD VDD P_18 W=10u L=1u m=1
MM3 Vx Vx VDD VDD P_18 W=10u L=1u m=1
MM2 Vout Vin2 Vp GND N_18 W=4u L=1u m=1
MM1 Vx Vin1 Vp GND N_18 W=4u L=1u m=1
.ENDS

