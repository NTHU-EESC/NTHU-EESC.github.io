************************************************************************
* Library Name: Lab1
* Cell Name:    FF
* View Name:    schematic
************************************************************************

.subckt FF vdd vss PRE CLK D CLR Q Qt
.param Wn13=3u Ln1=0.18u Wp13=2u Lp1=0.18u m1=1
.param Wn12=2u Wp12=2u

M1n11 out1 PRE n11 n11 n_18 W=Wn13 L=Ln1 m=m1
M1n12 n11 out4 n12 n12 n_18 W=Wn13 L=Ln1 m=m1
M1n13 n12 out2 vss vss n_18 W=Wn13 L=Ln1 m=m1
M1p11 out1 PRE vdd vdd p_18 W=Wp13 L=Lp1 m=m1
M1p12 out1 out4 vdd vdd p_18 W=Wp13 L=Lp1 m=m1
M1p13 out1 out2 vdd vdd p_18 W=Wp13 L=Lp1 m=m1

M1n21 out2 out1 n21 n21 n_18 W=Wn13 L=Ln1 m=m1
M1n22 n21 CLR n22 n22 n_18 W=Wn13 L=Ln1 m=m1
M1n23 n22 CLK vss vss n_18 W=Wn13 L=Ln1 m=m1
M1p21 out2 out1 vdd vdd p_18 W=Wp13 L=Lp1 m=m1
M1p22 out2 CLR vdd vdd p_18 W=Wp13 L=Lp1 m=m1
M1p23 out2 CLK vdd vdd p_18 W=Wp13 L=Lp1 m=m1

M1n31 out3 out2 n31 n31 n_18 W=Wn13 L=Ln1 m=m1
M1n32 n31 CLK n32 n32 n_18 W=Wn13 L=Ln1 m=m1
M1n33 n32 out4 vss vss n_18 W=Wn13 L=Ln1 m=m1
M1p31 out3 out2 vdd vdd p_18 W=Wp13 L=Lp1 m=m1
M1p32 out3 CLK vdd vdd p_18 W=Wp13 L=Lp1 m=m1
M1p33 out3 out4 vdd vdd p_18 W=Wp13 L=Lp1 m=m1

M1n41 out4 out3 n41 n41 n_18 W=Wn12 L=Ln1 m=m1
M1n42 n41 D vss vss n_18 W=Wn12 L=Ln1 m=m1
M1p41 out4 out3 vdd vdd p_18 W=Wp12 L=Lp1 m=m1
M1p42 out4 D vdd vdd p_18 W=Wp12 L=Lp1 m=m1

M1n51 Q PRE n51 n51 n_18 W=Wn13 L=Ln1 m=m1
M1n52 n51 out2 n52 n52 n_18 W=Wn13 L=Ln1 m=m1
M1n53 n52 Qt vss vss n_18 W=Wn13 L=Ln1 m=m1
M1p51 Q PRE vdd vdd p_18 W=Wp13 L=Lp1 m=m1
M1p52 Q out2 vdd vdd p_18 W=Wp13 L=Lp1 m=m1
M1p53 Q Qt vdd vdd p_18 W=Wp13 L=Lp1 m=m1

M1n61 Qt Q n61 n61 n_18 W=Wn13 L=Ln1 m=m1
M1n62 n61 out3 n62 n62 n_18 W=Wn13 L=Ln1 m=m1
M1n63 n62 CLR vss vss n_18 W=Wn13 L=Ln1 m=m1
M1p61 Qt Q vdd vdd p_18 W=Wp13 L=Lp1 m=m1
M1p62 Qt out3 vdd vdd p_18 W=Wp13 L=Lp1 m=m1
M1p63 Qt CLR vdd vdd p_18 W=Wp13 L=Lp1 m=m1

.ends


