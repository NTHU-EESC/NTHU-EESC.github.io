************************************************************************
* auCdl Netlist:
* 
* Library Name:  Hw2_1_a
* Top Cell Name: common_source
* View Name:     schematic
* Netlisted on:  Apr  1 19:49:28 2015
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: Hw2_1_a
* Cell Name:    common_source
* View Name:    schematic
************************************************************************

.SUBCKT common_source GND Vin Vout
*.PININFO GND:I Vin:I Vout:O
MM1 Vout Vin GND GND N_18 W=7.5u L=3u m=1
.ENDS

