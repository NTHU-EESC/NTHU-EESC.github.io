************************************************************************
* Library Name: 
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.subckt NAND2 vdd vss in1 in2 out
.param Wn13=3u Ln1=0.18u Wp13=2u Lp1=0.18u m1=1
.param Wn12=2u Wp12=2u

Mn1 out in1  n1  n1 n_18 W=2u L=2u m=m1
Mn2  n1 in2 vss vss n_18 W=2u L=2u m=m1
Mp1 out in1 vdd vdd p_18 W=2u L=2u m=m1
Mp2 out in2 vdd vdd p_18 W=2u L=2u m=m1

.ends


