* File: inv_chain2.pex.spi
* Created: Fri Dec  7 14:20:57 2018
* Program "Calibre xRC"
* Version "v2016.4_15.11"
* 
.include "inv_chain2.pex.spi.pex"
.subckt inv_chain2  VSS VDD OUT1 OUT2 OUT3 OUT4 OUT5 OUT9 OUT6 OUT7 OUT8
* 
* OUT8	OUT8
* OUT7	OUT7
* OUT6	OUT6
* OUT9	OUT9
* OUT5	OUT5
* OUT4	OUT4
* OUT3	OUT3
* OUT2	OUT2
* OUT1	OUT1
* VDD	VDD
* VSS	VSS
Mn1 N_OUT1_Mn1_d N_OUT9_Mn1_g N_VSS_Mn1_s N_VSS_Mn7@1159_b N_18 L=1.8e-07
+ W=5e-07 AD=2.955e-13 AS=2.995e-13 PD=1.682e-06 PS=1.698e-06
Mn2 N_OUT2_Mn2_d N_OUT1_Mn2_g N_VSS_Mn2_s N_VSS_Mn7@1159_b N_18 L=1.8e-07
+ W=5e-07 AD=1.325e-13 AS=2.995e-13 PD=5.3e-07 PS=1.698e-06
Mn2@3 N_OUT2_Mn2@3_d N_OUT1_Mn2@3_g N_VSS_Mn2@3_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.3125e-13 PD=5.3e-07 PS=5.25e-07
Mn2@2 N_OUT2_Mn2@2_d N_OUT1_Mn2@2_g N_VSS_Mn2@2_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=2.955e-13 AS=1.3125e-13 PD=1.682e-06 PS=5.25e-07
Mn3 N_OUT3_Mn3_d N_OUT2_Mn3_g N_VSS_Mn3_s N_VSS_Mn7@1159_b N_18 L=1.8e-07
+ W=5e-07 AD=1.325e-13 AS=2.995e-13 PD=5.3e-07 PS=1.698e-06
Mn3@11 N_OUT3_Mn3@11_d N_OUT2_Mn3@11_g N_VSS_Mn3@11_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn3@10 N_OUT3_Mn3@10_d N_OUT2_Mn3@10_g N_VSS_Mn3@10_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn3@9 N_OUT3_Mn3@9_d N_OUT2_Mn3@9_g N_VSS_Mn3@9_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn3@8 N_OUT3_Mn3@8_d N_OUT2_Mn3@8_g N_VSS_Mn3@8_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn3@7 N_OUT3_Mn3@7_d N_OUT2_Mn3@7_g N_VSS_Mn3@7_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn3@6 N_OUT3_Mn3@6_d N_OUT2_Mn3@6_g N_VSS_Mn3@6_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn3@5 N_OUT3_Mn3@5_d N_OUT2_Mn3@5_g N_VSS_Mn3@5_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn3@4 N_OUT3_Mn3@4_d N_OUT2_Mn3@4_g N_VSS_Mn3@4_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn3@3 N_OUT3_Mn3@3_d N_OUT2_Mn3@3_g N_VSS_Mn3@3_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn3@2 N_OUT3_Mn3@2_d N_OUT2_Mn3@2_g N_VSS_Mn3@2_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=2.955e-13 AS=1.4125e-13 PD=1.682e-06 PS=5.65e-07
Mn4 N_OUT4_Mn4_d N_OUT3_Mn4_g N_VSS_Mn4_s N_VSS_Mn7@1159_b N_18 L=1.8e-07
+ W=5e-07 AD=1.325e-13 AS=2.995e-13 PD=5.3e-07 PS=1.698e-06
Mn4@34 N_OUT4_Mn4@34_d N_OUT3_Mn4@34_g N_VSS_Mn4@34_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@33 N_OUT4_Mn4@33_d N_OUT3_Mn4@33_g N_VSS_Mn4@33_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@32 N_OUT4_Mn4@32_d N_OUT3_Mn4@32_g N_VSS_Mn4@32_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@31 N_OUT4_Mn4@31_d N_OUT3_Mn4@31_g N_VSS_Mn4@31_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@30 N_OUT4_Mn4@30_d N_OUT3_Mn4@30_g N_VSS_Mn4@30_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@29 N_OUT4_Mn4@29_d N_OUT3_Mn4@29_g N_VSS_Mn4@29_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@28 N_OUT4_Mn4@28_d N_OUT3_Mn4@28_g N_VSS_Mn4@28_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@27 N_OUT4_Mn4@27_d N_OUT3_Mn4@27_g N_VSS_Mn4@27_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@26 N_OUT4_Mn4@26_d N_OUT3_Mn4@26_g N_VSS_Mn4@26_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@25 N_OUT4_Mn4@25_d N_OUT3_Mn4@25_g N_VSS_Mn4@25_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@24 N_OUT4_Mn4@24_d N_OUT3_Mn4@24_g N_VSS_Mn4@24_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@23 N_OUT4_Mn4@23_d N_OUT3_Mn4@23_g N_VSS_Mn4@23_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@22 N_OUT4_Mn4@22_d N_OUT3_Mn4@22_g N_VSS_Mn4@22_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@21 N_OUT4_Mn4@21_d N_OUT3_Mn4@21_g N_VSS_Mn4@21_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@20 N_OUT4_Mn4@20_d N_OUT3_Mn4@20_g N_VSS_Mn4@20_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@19 N_OUT4_Mn4@19_d N_OUT3_Mn4@19_g N_VSS_Mn4@19_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@18 N_OUT4_Mn4@18_d N_OUT3_Mn4@18_g N_VSS_Mn4@18_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@17 N_OUT4_Mn4@17_d N_OUT3_Mn4@17_g N_VSS_Mn4@17_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@16 N_OUT4_Mn4@16_d N_OUT3_Mn4@16_g N_VSS_Mn4@16_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@15 N_OUT4_Mn4@15_d N_OUT3_Mn4@15_g N_VSS_Mn4@15_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@14 N_OUT4_Mn4@14_d N_OUT3_Mn4@14_g N_VSS_Mn4@14_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@13 N_OUT4_Mn4@13_d N_OUT3_Mn4@13_g N_VSS_Mn4@13_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@12 N_OUT4_Mn4@12_d N_OUT3_Mn4@12_g N_VSS_Mn4@12_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@11 N_OUT4_Mn4@11_d N_OUT3_Mn4@11_g N_VSS_Mn4@11_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@10 N_OUT4_Mn4@10_d N_OUT3_Mn4@10_g N_VSS_Mn4@10_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@9 N_OUT4_Mn4@9_d N_OUT3_Mn4@9_g N_VSS_Mn4@9_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@8 N_OUT4_Mn4@8_d N_OUT3_Mn4@8_g N_VSS_Mn4@8_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@7 N_OUT4_Mn4@7_d N_OUT3_Mn4@7_g N_VSS_Mn4@7_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@6 N_OUT4_Mn4@6_d N_OUT3_Mn4@6_g N_VSS_Mn4@6_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@5 N_OUT4_Mn4@5_d N_OUT3_Mn4@5_g N_VSS_Mn4@5_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn4@4 N_OUT4_Mn4@4_d N_OUT3_Mn4@4_g N_VSS_Mn4@4_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.275e-13 PD=5.3e-07 PS=5.1e-07
Mn4@3 N_OUT4_Mn4@3_d N_OUT3_Mn4@3_g N_VSS_Mn4@3_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.4375e-13 AS=1.275e-13 PD=5.75e-07 PS=5.1e-07
Mn4@2 N_OUT4_Mn4@2_d N_OUT3_Mn4@2_g N_VSS_Mn4@2_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.4375e-13 AS=3.005e-13 PD=5.75e-07 PS=1.702e-06
Mn5 N_OUT5_Mn5_d N_OUT4_Mn5_g N_VSS_Mn5_s N_VSS_Mn7@1159_b N_18 L=1.8e-07
+ W=5e-07 AD=1.325e-13 AS=2.995e-13 PD=5.3e-07 PS=1.698e-06
Mn5@111 N_OUT5_Mn5@111_d N_OUT4_Mn5@111_g N_VSS_Mn5@111_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@110 N_OUT5_Mn5@110_d N_OUT4_Mn5@110_g N_VSS_Mn5@110_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@109 N_OUT5_Mn5@109_d N_OUT4_Mn5@109_g N_VSS_Mn5@109_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@108 N_OUT5_Mn5@108_d N_OUT4_Mn5@108_g N_VSS_Mn5@108_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@107 N_OUT5_Mn5@107_d N_OUT4_Mn5@107_g N_VSS_Mn5@107_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@106 N_OUT5_Mn5@106_d N_OUT4_Mn5@106_g N_VSS_Mn5@106_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=2.955e-13 AS=1.4125e-13 PD=1.682e-06 PS=5.65e-07
Mn6 N_OUT6_Mn6_d N_OUT5_Mn6_g N_VSS_Mn6_s N_VSS_Mn7@1159_b N_18 L=1.8e-07
+ W=5e-07 AD=1.325e-13 AS=2.995e-13 PD=5.3e-07 PS=1.698e-06
Mn9 N_OUT9_Mn9_d N_OUT8_Mn9_g N_VSS_Mn9_s N_VSS_Mn7@1159_b N_18 L=1.8e-07
+ W=1.1e-06 AD=6.501e-13 AS=3.1075e-13 PD=2.282e-06 PS=5.65e-07
Mn6@359 N_OUT6_Mn6@359_d N_OUT5_Mn6@359_g N_VSS_Mn6@359_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@358 N_OUT6_Mn6@358_d N_OUT5_Mn6@358_g N_VSS_Mn6@358_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@357 N_OUT6_Mn6@357_d N_OUT5_Mn6@357_g N_VSS_Mn6@357_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@356 N_OUT6_Mn6@356_d N_OUT5_Mn6@356_g N_VSS_Mn6@356_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@355 N_OUT6_Mn6@355_d N_OUT5_Mn6@355_g N_VSS_Mn6@355_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@354 N_OUT6_Mn6@354_d N_OUT5_Mn6@354_g N_VSS_Mn6@354_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@353 N_OUT6_Mn6@353_d N_OUT5_Mn6@353_g N_VSS_Mn6@353_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@352 N_OUT6_Mn6@352_d N_OUT5_Mn6@352_g N_VSS_Mn6@352_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@351 N_OUT6_Mn6@351_d N_OUT5_Mn6@351_g N_VSS_Mn6@351_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@350 N_OUT6_Mn6@350_d N_OUT5_Mn6@350_g N_VSS_Mn6@350_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@349 N_OUT6_Mn6@349_d N_OUT5_Mn6@349_g N_VSS_Mn6@349_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@348 N_OUT6_Mn6@348_d N_OUT5_Mn6@348_g N_VSS_Mn6@348_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@347 N_OUT6_Mn6@347_d N_OUT5_Mn6@347_g N_VSS_Mn6@347_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@346 N_OUT6_Mn6@346_d N_OUT5_Mn6@346_g N_VSS_Mn6@346_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@345 N_OUT6_Mn6@345_d N_OUT5_Mn6@345_g N_VSS_Mn6@345_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@344 N_OUT6_Mn6@344_d N_OUT5_Mn6@344_g N_VSS_Mn6@344_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@343 N_OUT6_Mn6@343_d N_OUT5_Mn6@343_g N_VSS_Mn6@343_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@342 N_OUT6_Mn6@342_d N_OUT5_Mn6@342_g N_VSS_Mn6@342_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@341 N_OUT6_Mn6@341_d N_OUT5_Mn6@341_g N_VSS_Mn6@341_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@340 N_OUT6_Mn6@340_d N_OUT5_Mn6@340_g N_VSS_Mn6@340_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@339 N_OUT6_Mn6@339_d N_OUT5_Mn6@339_g N_VSS_Mn6@339_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@338 N_OUT6_Mn6@338_d N_OUT5_Mn6@338_g N_VSS_Mn6@338_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@337 N_OUT6_Mn6@337_d N_OUT5_Mn6@337_g N_VSS_Mn6@337_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@336 N_OUT6_Mn6@336_d N_OUT5_Mn6@336_g N_VSS_Mn6@336_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@335 N_OUT6_Mn6@335_d N_OUT5_Mn6@335_g N_VSS_Mn6@335_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@334 N_OUT6_Mn6@334_d N_OUT5_Mn6@334_g N_VSS_Mn6@334_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@333 N_OUT6_Mn6@333_d N_OUT5_Mn6@333_g N_VSS_Mn6@333_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@332 N_OUT6_Mn6@332_d N_OUT5_Mn6@332_g N_VSS_Mn6@332_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@331 N_OUT6_Mn6@331_d N_OUT5_Mn6@331_g N_VSS_Mn6@331_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@330 N_OUT6_Mn6@330_d N_OUT5_Mn6@330_g N_VSS_Mn6@330_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@329 N_OUT6_Mn6@329_d N_OUT5_Mn6@329_g N_VSS_Mn6@329_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@328 N_OUT6_Mn6@328_d N_OUT5_Mn6@328_g N_VSS_Mn6@328_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@327 N_OUT6_Mn6@327_d N_OUT5_Mn6@327_g N_VSS_Mn6@327_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@326 N_OUT6_Mn6@326_d N_OUT5_Mn6@326_g N_VSS_Mn6@326_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@325 N_OUT6_Mn6@325_d N_OUT5_Mn6@325_g N_VSS_Mn6@325_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@324 N_OUT6_Mn6@324_d N_OUT5_Mn6@324_g N_VSS_Mn6@324_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@323 N_OUT6_Mn6@323_d N_OUT5_Mn6@323_g N_VSS_Mn6@323_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@322 N_OUT6_Mn6@322_d N_OUT5_Mn6@322_g N_VSS_Mn6@322_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@321 N_OUT6_Mn6@321_d N_OUT5_Mn6@321_g N_VSS_Mn6@321_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@320 N_OUT6_Mn6@320_d N_OUT5_Mn6@320_g N_VSS_Mn6@320_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@319 N_OUT6_Mn6@319_d N_OUT5_Mn6@319_g N_VSS_Mn6@319_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@318 N_OUT6_Mn6@318_d N_OUT5_Mn6@318_g N_VSS_Mn6@318_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@317 N_OUT6_Mn6@317_d N_OUT5_Mn6@317_g N_VSS_Mn6@317_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@316 N_OUT6_Mn6@316_d N_OUT5_Mn6@316_g N_VSS_Mn6@316_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@315 N_OUT6_Mn6@315_d N_OUT5_Mn6@315_g N_VSS_Mn6@315_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@314 N_OUT6_Mn6@314_d N_OUT5_Mn6@314_g N_VSS_Mn6@314_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@313 N_OUT6_Mn6@313_d N_OUT5_Mn6@313_g N_VSS_Mn6@313_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@312 N_OUT6_Mn6@312_d N_OUT5_Mn6@312_g N_VSS_Mn6@312_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@311 N_OUT6_Mn6@311_d N_OUT5_Mn6@311_g N_VSS_Mn6@311_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@310 N_OUT6_Mn6@310_d N_OUT5_Mn6@310_g N_VSS_Mn6@310_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@309 N_OUT6_Mn6@309_d N_OUT5_Mn6@309_g N_VSS_Mn6@309_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@308 N_OUT6_Mn6@308_d N_OUT5_Mn6@308_g N_VSS_Mn6@308_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@307 N_OUT6_Mn6@307_d N_OUT5_Mn6@307_g N_VSS_Mn6@307_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@306 N_OUT6_Mn6@306_d N_OUT5_Mn6@306_g N_VSS_Mn6@306_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@305 N_OUT6_Mn6@305_d N_OUT5_Mn6@305_g N_VSS_Mn6@305_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@304 N_OUT6_Mn6@304_d N_OUT5_Mn6@304_g N_VSS_Mn6@304_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@303 N_OUT6_Mn6@303_d N_OUT5_Mn6@303_g N_VSS_Mn6@303_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@302 N_OUT6_Mn6@302_d N_OUT5_Mn6@302_g N_VSS_Mn6@302_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@301 N_OUT6_Mn6@301_d N_OUT5_Mn6@301_g N_VSS_Mn6@301_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@300 N_OUT6_Mn6@300_d N_OUT5_Mn6@300_g N_VSS_Mn6@300_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@299 N_OUT6_Mn6@299_d N_OUT5_Mn6@299_g N_VSS_Mn6@299_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@298 N_OUT6_Mn6@298_d N_OUT5_Mn6@298_g N_VSS_Mn6@298_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@297 N_OUT6_Mn6@297_d N_OUT5_Mn6@297_g N_VSS_Mn6@297_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@296 N_OUT6_Mn6@296_d N_OUT5_Mn6@296_g N_VSS_Mn6@296_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@295 N_OUT6_Mn6@295_d N_OUT5_Mn6@295_g N_VSS_Mn6@295_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@294 N_OUT6_Mn6@294_d N_OUT5_Mn6@294_g N_VSS_Mn6@294_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@293 N_OUT6_Mn6@293_d N_OUT5_Mn6@293_g N_VSS_Mn6@293_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@292 N_OUT6_Mn6@292_d N_OUT5_Mn6@292_g N_VSS_Mn6@292_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@291 N_OUT6_Mn6@291_d N_OUT5_Mn6@291_g N_VSS_Mn6@291_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@290 N_OUT6_Mn6@290_d N_OUT5_Mn6@290_g N_VSS_Mn6@290_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@289 N_OUT6_Mn6@289_d N_OUT5_Mn6@289_g N_VSS_Mn6@289_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@288 N_OUT6_Mn6@288_d N_OUT5_Mn6@288_g N_VSS_Mn6@288_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@287 N_OUT6_Mn6@287_d N_OUT5_Mn6@287_g N_VSS_Mn6@287_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@286 N_OUT6_Mn6@286_d N_OUT5_Mn6@286_g N_VSS_Mn6@286_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@285 N_OUT6_Mn6@285_d N_OUT5_Mn6@285_g N_VSS_Mn6@285_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@284 N_OUT6_Mn6@284_d N_OUT5_Mn6@284_g N_VSS_Mn6@284_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@283 N_OUT6_Mn6@283_d N_OUT5_Mn6@283_g N_VSS_Mn6@283_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@282 N_OUT6_Mn6@282_d N_OUT5_Mn6@282_g N_VSS_Mn6@282_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@281 N_OUT6_Mn6@281_d N_OUT5_Mn6@281_g N_VSS_Mn6@281_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@280 N_OUT6_Mn6@280_d N_OUT5_Mn6@280_g N_VSS_Mn6@280_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@279 N_OUT6_Mn6@279_d N_OUT5_Mn6@279_g N_VSS_Mn6@279_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@278 N_OUT6_Mn6@278_d N_OUT5_Mn6@278_g N_VSS_Mn6@278_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@277 N_OUT6_Mn6@277_d N_OUT5_Mn6@277_g N_VSS_Mn6@277_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@276 N_OUT6_Mn6@276_d N_OUT5_Mn6@276_g N_VSS_Mn6@276_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@275 N_OUT6_Mn6@275_d N_OUT5_Mn6@275_g N_VSS_Mn6@275_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@274 N_OUT6_Mn6@274_d N_OUT5_Mn6@274_g N_VSS_Mn6@274_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@273 N_OUT6_Mn6@273_d N_OUT5_Mn6@273_g N_VSS_Mn6@273_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@272 N_OUT6_Mn6@272_d N_OUT5_Mn6@272_g N_VSS_Mn6@272_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@271 N_OUT6_Mn6@271_d N_OUT5_Mn6@271_g N_VSS_Mn6@271_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@270 N_OUT6_Mn6@270_d N_OUT5_Mn6@270_g N_VSS_Mn6@270_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@269 N_OUT6_Mn6@269_d N_OUT5_Mn6@269_g N_VSS_Mn6@269_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@268 N_OUT6_Mn6@268_d N_OUT5_Mn6@268_g N_VSS_Mn6@268_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@267 N_OUT6_Mn6@267_d N_OUT5_Mn6@267_g N_VSS_Mn6@267_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@266 N_OUT6_Mn6@266_d N_OUT5_Mn6@266_g N_VSS_Mn6@266_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@265 N_OUT6_Mn6@265_d N_OUT5_Mn6@265_g N_VSS_Mn6@265_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@264 N_OUT6_Mn6@264_d N_OUT5_Mn6@264_g N_VSS_Mn6@264_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@263 N_OUT6_Mn6@263_d N_OUT5_Mn6@263_g N_VSS_Mn6@263_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@262 N_OUT6_Mn6@262_d N_OUT5_Mn6@262_g N_VSS_Mn6@262_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@261 N_OUT6_Mn6@261_d N_OUT5_Mn6@261_g N_VSS_Mn6@261_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@260 N_OUT6_Mn6@260_d N_OUT5_Mn6@260_g N_VSS_Mn6@260_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@259 N_OUT6_Mn6@259_d N_OUT5_Mn6@259_g N_VSS_Mn6@259_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@258 N_OUT6_Mn6@258_d N_OUT5_Mn6@258_g N_VSS_Mn6@258_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@257 N_OUT6_Mn6@257_d N_OUT5_Mn6@257_g N_VSS_Mn6@257_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@256 N_OUT6_Mn6@256_d N_OUT5_Mn6@256_g N_VSS_Mn6@256_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@255 N_OUT6_Mn6@255_d N_OUT5_Mn6@255_g N_VSS_Mn6@255_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@254 N_OUT6_Mn6@254_d N_OUT5_Mn6@254_g N_VSS_Mn6@254_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@253 N_OUT6_Mn6@253_d N_OUT5_Mn6@253_g N_VSS_Mn6@253_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@252 N_OUT6_Mn6@252_d N_OUT5_Mn6@252_g N_VSS_Mn6@252_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@251 N_OUT6_Mn6@251_d N_OUT5_Mn6@251_g N_VSS_Mn6@251_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@250 N_OUT6_Mn6@250_d N_OUT5_Mn6@250_g N_VSS_Mn6@250_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@249 N_OUT6_Mn6@249_d N_OUT5_Mn6@249_g N_VSS_Mn6@249_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@248 N_OUT6_Mn6@248_d N_OUT5_Mn6@248_g N_VSS_Mn6@248_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@247 N_OUT6_Mn6@247_d N_OUT5_Mn6@247_g N_VSS_Mn6@247_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@246 N_OUT6_Mn6@246_d N_OUT5_Mn6@246_g N_VSS_Mn6@246_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@245 N_OUT6_Mn6@245_d N_OUT5_Mn6@245_g N_VSS_Mn6@245_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@244 N_OUT6_Mn6@244_d N_OUT5_Mn6@244_g N_VSS_Mn6@244_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@243 N_OUT6_Mn6@243_d N_OUT5_Mn6@243_g N_VSS_Mn6@243_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@242 N_OUT6_Mn6@242_d N_OUT5_Mn6@242_g N_VSS_Mn6@242_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@241 N_OUT6_Mn6@241_d N_OUT5_Mn6@241_g N_VSS_Mn6@241_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@240 N_OUT6_Mn6@240_d N_OUT5_Mn6@240_g N_VSS_Mn6@240_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@239 N_OUT6_Mn6@239_d N_OUT5_Mn6@239_g N_VSS_Mn6@239_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@238 N_OUT6_Mn6@238_d N_OUT5_Mn6@238_g N_VSS_Mn6@238_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@237 N_OUT6_Mn6@237_d N_OUT5_Mn6@237_g N_VSS_Mn6@237_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@236 N_OUT6_Mn6@236_d N_OUT5_Mn6@236_g N_VSS_Mn6@236_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@235 N_OUT6_Mn6@235_d N_OUT5_Mn6@235_g N_VSS_Mn6@235_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@234 N_OUT6_Mn6@234_d N_OUT5_Mn6@234_g N_VSS_Mn6@234_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@233 N_OUT6_Mn6@233_d N_OUT5_Mn6@233_g N_VSS_Mn6@233_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@232 N_OUT6_Mn6@232_d N_OUT5_Mn6@232_g N_VSS_Mn6@232_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@231 N_OUT6_Mn6@231_d N_OUT5_Mn6@231_g N_VSS_Mn6@231_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@230 N_OUT6_Mn6@230_d N_OUT5_Mn6@230_g N_VSS_Mn6@230_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@229 N_OUT6_Mn6@229_d N_OUT5_Mn6@229_g N_VSS_Mn6@229_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@228 N_OUT6_Mn6@228_d N_OUT5_Mn6@228_g N_VSS_Mn6@228_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@227 N_OUT6_Mn6@227_d N_OUT5_Mn6@227_g N_VSS_Mn6@227_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@226 N_OUT6_Mn6@226_d N_OUT5_Mn6@226_g N_VSS_Mn6@226_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@225 N_OUT6_Mn6@225_d N_OUT5_Mn6@225_g N_VSS_Mn6@225_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@224 N_OUT6_Mn6@224_d N_OUT5_Mn6@224_g N_VSS_Mn6@224_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@223 N_OUT6_Mn6@223_d N_OUT5_Mn6@223_g N_VSS_Mn6@223_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@222 N_OUT6_Mn6@222_d N_OUT5_Mn6@222_g N_VSS_Mn6@222_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@221 N_OUT6_Mn6@221_d N_OUT5_Mn6@221_g N_VSS_Mn6@221_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@220 N_OUT6_Mn6@220_d N_OUT5_Mn6@220_g N_VSS_Mn6@220_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@219 N_OUT6_Mn6@219_d N_OUT5_Mn6@219_g N_VSS_Mn6@219_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@218 N_OUT6_Mn6@218_d N_OUT5_Mn6@218_g N_VSS_Mn6@218_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@217 N_OUT6_Mn6@217_d N_OUT5_Mn6@217_g N_VSS_Mn6@217_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@216 N_OUT6_Mn6@216_d N_OUT5_Mn6@216_g N_VSS_Mn6@216_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@215 N_OUT6_Mn6@215_d N_OUT5_Mn6@215_g N_VSS_Mn6@215_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@214 N_OUT6_Mn6@214_d N_OUT5_Mn6@214_g N_VSS_Mn6@214_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@213 N_OUT6_Mn6@213_d N_OUT5_Mn6@213_g N_VSS_Mn6@213_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@212 N_OUT6_Mn6@212_d N_OUT5_Mn6@212_g N_VSS_Mn6@212_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@211 N_OUT6_Mn6@211_d N_OUT5_Mn6@211_g N_VSS_Mn6@211_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@210 N_OUT6_Mn6@210_d N_OUT5_Mn6@210_g N_VSS_Mn6@210_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@209 N_OUT6_Mn6@209_d N_OUT5_Mn6@209_g N_VSS_Mn6@209_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@208 N_OUT6_Mn6@208_d N_OUT5_Mn6@208_g N_VSS_Mn6@208_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@207 N_OUT6_Mn6@207_d N_OUT5_Mn6@207_g N_VSS_Mn6@207_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@206 N_OUT6_Mn6@206_d N_OUT5_Mn6@206_g N_VSS_Mn6@206_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@205 N_OUT6_Mn6@205_d N_OUT5_Mn6@205_g N_VSS_Mn6@205_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@204 N_OUT6_Mn6@204_d N_OUT5_Mn6@204_g N_VSS_Mn6@204_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@203 N_OUT6_Mn6@203_d N_OUT5_Mn6@203_g N_VSS_Mn6@203_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@202 N_OUT6_Mn6@202_d N_OUT5_Mn6@202_g N_VSS_Mn6@202_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@201 N_OUT6_Mn6@201_d N_OUT5_Mn6@201_g N_VSS_Mn6@201_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@200 N_OUT6_Mn6@200_d N_OUT5_Mn6@200_g N_VSS_Mn6@200_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@199 N_OUT6_Mn6@199_d N_OUT5_Mn6@199_g N_VSS_Mn6@199_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@198 N_OUT6_Mn6@198_d N_OUT5_Mn6@198_g N_VSS_Mn6@198_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@197 N_OUT6_Mn6@197_d N_OUT5_Mn6@197_g N_VSS_Mn6@197_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@196 N_OUT6_Mn6@196_d N_OUT5_Mn6@196_g N_VSS_Mn6@196_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@195 N_OUT6_Mn6@195_d N_OUT5_Mn6@195_g N_VSS_Mn6@195_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@194 N_OUT6_Mn6@194_d N_OUT5_Mn6@194_g N_VSS_Mn6@194_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@193 N_OUT6_Mn6@193_d N_OUT5_Mn6@193_g N_VSS_Mn6@193_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@192 N_OUT6_Mn6@192_d N_OUT5_Mn6@192_g N_VSS_Mn6@192_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@191 N_OUT6_Mn6@191_d N_OUT5_Mn6@191_g N_VSS_Mn6@191_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@190 N_OUT6_Mn6@190_d N_OUT5_Mn6@190_g N_VSS_Mn6@190_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@189 N_OUT6_Mn6@189_d N_OUT5_Mn6@189_g N_VSS_Mn6@189_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@188 N_OUT6_Mn6@188_d N_OUT5_Mn6@188_g N_VSS_Mn6@188_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@187 N_OUT6_Mn6@187_d N_OUT5_Mn6@187_g N_VSS_Mn6@187_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@186 N_OUT6_Mn6@186_d N_OUT5_Mn6@186_g N_VSS_Mn6@186_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@185 N_OUT6_Mn6@185_d N_OUT5_Mn6@185_g N_VSS_Mn6@185_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@184 N_OUT6_Mn6@184_d N_OUT5_Mn6@184_g N_VSS_Mn6@184_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@183 N_OUT6_Mn6@183_d N_OUT5_Mn6@183_g N_VSS_Mn6@183_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@182 N_OUT6_Mn6@182_d N_OUT5_Mn6@182_g N_VSS_Mn6@182_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@181 N_OUT6_Mn6@181_d N_OUT5_Mn6@181_g N_VSS_Mn6@181_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@180 N_OUT6_Mn6@180_d N_OUT5_Mn6@180_g N_VSS_Mn6@180_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@179 N_OUT6_Mn6@179_d N_OUT5_Mn6@179_g N_VSS_Mn6@179_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@178 N_OUT6_Mn6@178_d N_OUT5_Mn6@178_g N_VSS_Mn6@178_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@177 N_OUT6_Mn6@177_d N_OUT5_Mn6@177_g N_VSS_Mn6@177_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@176 N_OUT6_Mn6@176_d N_OUT5_Mn6@176_g N_VSS_Mn6@176_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@175 N_OUT6_Mn6@175_d N_OUT5_Mn6@175_g N_VSS_Mn6@175_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@174 N_OUT6_Mn6@174_d N_OUT5_Mn6@174_g N_VSS_Mn6@174_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@173 N_OUT6_Mn6@173_d N_OUT5_Mn6@173_g N_VSS_Mn6@173_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@172 N_OUT6_Mn6@172_d N_OUT5_Mn6@172_g N_VSS_Mn6@172_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@171 N_OUT6_Mn6@171_d N_OUT5_Mn6@171_g N_VSS_Mn6@171_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@170 N_OUT6_Mn6@170_d N_OUT5_Mn6@170_g N_VSS_Mn6@170_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@169 N_OUT6_Mn6@169_d N_OUT5_Mn6@169_g N_VSS_Mn6@169_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@168 N_OUT6_Mn6@168_d N_OUT5_Mn6@168_g N_VSS_Mn6@168_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@167 N_OUT6_Mn6@167_d N_OUT5_Mn6@167_g N_VSS_Mn6@167_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@166 N_OUT6_Mn6@166_d N_OUT5_Mn6@166_g N_VSS_Mn6@166_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@165 N_OUT6_Mn6@165_d N_OUT5_Mn6@165_g N_VSS_Mn6@165_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@164 N_OUT6_Mn6@164_d N_OUT5_Mn6@164_g N_VSS_Mn6@164_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@163 N_OUT6_Mn6@163_d N_OUT5_Mn6@163_g N_VSS_Mn6@163_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@162 N_OUT6_Mn6@162_d N_OUT5_Mn6@162_g N_VSS_Mn6@162_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@161 N_OUT6_Mn6@161_d N_OUT5_Mn6@161_g N_VSS_Mn6@161_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@160 N_OUT6_Mn6@160_d N_OUT5_Mn6@160_g N_VSS_Mn6@160_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@159 N_OUT6_Mn6@159_d N_OUT5_Mn6@159_g N_VSS_Mn6@159_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@158 N_OUT6_Mn6@158_d N_OUT5_Mn6@158_g N_VSS_Mn6@158_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@157 N_OUT6_Mn6@157_d N_OUT5_Mn6@157_g N_VSS_Mn6@157_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@156 N_OUT6_Mn6@156_d N_OUT5_Mn6@156_g N_VSS_Mn6@156_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@155 N_OUT6_Mn6@155_d N_OUT5_Mn6@155_g N_VSS_Mn6@155_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@154 N_OUT6_Mn6@154_d N_OUT5_Mn6@154_g N_VSS_Mn6@154_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@153 N_OUT6_Mn6@153_d N_OUT5_Mn6@153_g N_VSS_Mn6@153_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@152 N_OUT6_Mn6@152_d N_OUT5_Mn6@152_g N_VSS_Mn6@152_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@151 N_OUT6_Mn6@151_d N_OUT5_Mn6@151_g N_VSS_Mn6@151_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@150 N_OUT6_Mn6@150_d N_OUT5_Mn6@150_g N_VSS_Mn6@150_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@149 N_OUT6_Mn6@149_d N_OUT5_Mn6@149_g N_VSS_Mn6@149_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@148 N_OUT6_Mn6@148_d N_OUT5_Mn6@148_g N_VSS_Mn6@148_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@147 N_OUT6_Mn6@147_d N_OUT5_Mn6@147_g N_VSS_Mn6@147_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@146 N_OUT6_Mn6@146_d N_OUT5_Mn6@146_g N_VSS_Mn6@146_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@145 N_OUT6_Mn6@145_d N_OUT5_Mn6@145_g N_VSS_Mn6@145_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@144 N_OUT6_Mn6@144_d N_OUT5_Mn6@144_g N_VSS_Mn6@144_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@143 N_OUT6_Mn6@143_d N_OUT5_Mn6@143_g N_VSS_Mn6@143_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@142 N_OUT6_Mn6@142_d N_OUT5_Mn6@142_g N_VSS_Mn6@142_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@141 N_OUT6_Mn6@141_d N_OUT5_Mn6@141_g N_VSS_Mn6@141_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@140 N_OUT6_Mn6@140_d N_OUT5_Mn6@140_g N_VSS_Mn6@140_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@139 N_OUT6_Mn6@139_d N_OUT5_Mn6@139_g N_VSS_Mn6@139_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@138 N_OUT6_Mn6@138_d N_OUT5_Mn6@138_g N_VSS_Mn6@138_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@137 N_OUT6_Mn6@137_d N_OUT5_Mn6@137_g N_VSS_Mn6@137_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@136 N_OUT6_Mn6@136_d N_OUT5_Mn6@136_g N_VSS_Mn6@136_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@135 N_OUT6_Mn6@135_d N_OUT5_Mn6@135_g N_VSS_Mn6@135_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@134 N_OUT6_Mn6@134_d N_OUT5_Mn6@134_g N_VSS_Mn6@134_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@133 N_OUT6_Mn6@133_d N_OUT5_Mn6@133_g N_VSS_Mn6@133_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@132 N_OUT6_Mn6@132_d N_OUT5_Mn6@132_g N_VSS_Mn6@132_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@131 N_OUT6_Mn6@131_d N_OUT5_Mn6@131_g N_VSS_Mn6@131_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@130 N_OUT6_Mn6@130_d N_OUT5_Mn6@130_g N_VSS_Mn6@130_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@129 N_OUT6_Mn6@129_d N_OUT5_Mn6@129_g N_VSS_Mn6@129_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@128 N_OUT6_Mn6@128_d N_OUT5_Mn6@128_g N_VSS_Mn6@128_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@127 N_OUT6_Mn6@127_d N_OUT5_Mn6@127_g N_VSS_Mn6@127_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@126 N_OUT6_Mn6@126_d N_OUT5_Mn6@126_g N_VSS_Mn6@126_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@125 N_OUT6_Mn6@125_d N_OUT5_Mn6@125_g N_VSS_Mn6@125_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@124 N_OUT6_Mn6@124_d N_OUT5_Mn6@124_g N_VSS_Mn6@124_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@123 N_OUT6_Mn6@123_d N_OUT5_Mn6@123_g N_VSS_Mn6@123_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@122 N_OUT6_Mn6@122_d N_OUT5_Mn6@122_g N_VSS_Mn6@122_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@121 N_OUT6_Mn6@121_d N_OUT5_Mn6@121_g N_VSS_Mn6@121_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@120 N_OUT6_Mn6@120_d N_OUT5_Mn6@120_g N_VSS_Mn6@120_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@119 N_OUT6_Mn6@119_d N_OUT5_Mn6@119_g N_VSS_Mn6@119_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@118 N_OUT6_Mn6@118_d N_OUT5_Mn6@118_g N_VSS_Mn6@118_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@117 N_OUT6_Mn6@117_d N_OUT5_Mn6@117_g N_VSS_Mn6@117_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@116 N_OUT6_Mn6@116_d N_OUT5_Mn6@116_g N_VSS_Mn6@116_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@115 N_OUT6_Mn6@115_d N_OUT5_Mn6@115_g N_VSS_Mn6@115_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@114 N_OUT6_Mn6@114_d N_OUT5_Mn6@114_g N_VSS_Mn6@114_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@113 N_OUT6_Mn6@113_d N_OUT5_Mn6@113_g N_VSS_Mn6@113_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@112 N_OUT6_Mn6@112_d N_OUT5_Mn6@112_g N_VSS_Mn6@112_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@111 N_OUT6_Mn6@111_d N_OUT5_Mn6@111_g N_VSS_Mn6@111_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@110 N_OUT6_Mn6@110_d N_OUT5_Mn6@110_g N_VSS_Mn6@110_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@109 N_OUT6_Mn6@109_d N_OUT5_Mn6@109_g N_VSS_Mn6@109_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@108 N_OUT6_Mn6@108_d N_OUT5_Mn6@108_g N_VSS_Mn6@108_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@107 N_OUT6_Mn6@107_d N_OUT5_Mn6@107_g N_VSS_Mn6@107_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@106 N_OUT6_Mn6@106_d N_OUT5_Mn6@106_g N_VSS_Mn6@106_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@105 N_OUT6_Mn6@105_d N_OUT5_Mn6@105_g N_VSS_Mn6@105_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@104 N_OUT6_Mn6@104_d N_OUT5_Mn6@104_g N_VSS_Mn6@104_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@103 N_OUT6_Mn6@103_d N_OUT5_Mn6@103_g N_VSS_Mn6@103_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@102 N_OUT6_Mn6@102_d N_OUT5_Mn6@102_g N_VSS_Mn6@102_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@101 N_OUT6_Mn6@101_d N_OUT5_Mn6@101_g N_VSS_Mn6@101_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@100 N_OUT6_Mn6@100_d N_OUT5_Mn6@100_g N_VSS_Mn6@100_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@99 N_OUT6_Mn6@99_d N_OUT5_Mn6@99_g N_VSS_Mn6@99_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@98 N_OUT6_Mn6@98_d N_OUT5_Mn6@98_g N_VSS_Mn6@98_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@97 N_OUT6_Mn6@97_d N_OUT5_Mn6@97_g N_VSS_Mn6@97_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@96 N_OUT6_Mn6@96_d N_OUT5_Mn6@96_g N_VSS_Mn6@96_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@95 N_OUT6_Mn6@95_d N_OUT5_Mn6@95_g N_VSS_Mn6@95_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@94 N_OUT6_Mn6@94_d N_OUT5_Mn6@94_g N_VSS_Mn6@94_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@93 N_OUT6_Mn6@93_d N_OUT5_Mn6@93_g N_VSS_Mn6@93_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@92 N_OUT6_Mn6@92_d N_OUT5_Mn6@92_g N_VSS_Mn6@92_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@91 N_OUT6_Mn6@91_d N_OUT5_Mn6@91_g N_VSS_Mn6@91_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@90 N_OUT6_Mn6@90_d N_OUT5_Mn6@90_g N_VSS_Mn6@90_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@89 N_OUT6_Mn6@89_d N_OUT5_Mn6@89_g N_VSS_Mn6@89_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@88 N_OUT6_Mn6@88_d N_OUT5_Mn6@88_g N_VSS_Mn6@88_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@87 N_OUT6_Mn6@87_d N_OUT5_Mn6@87_g N_VSS_Mn6@87_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@86 N_OUT6_Mn6@86_d N_OUT5_Mn6@86_g N_VSS_Mn6@86_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@85 N_OUT6_Mn6@85_d N_OUT5_Mn6@85_g N_VSS_Mn6@85_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@84 N_OUT6_Mn6@84_d N_OUT5_Mn6@84_g N_VSS_Mn6@84_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@83 N_OUT6_Mn6@83_d N_OUT5_Mn6@83_g N_VSS_Mn6@83_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@82 N_OUT6_Mn6@82_d N_OUT5_Mn6@82_g N_VSS_Mn6@82_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@81 N_OUT6_Mn6@81_d N_OUT5_Mn6@81_g N_VSS_Mn6@81_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@80 N_OUT6_Mn6@80_d N_OUT5_Mn6@80_g N_VSS_Mn6@80_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@79 N_OUT6_Mn6@79_d N_OUT5_Mn6@79_g N_VSS_Mn6@79_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@78 N_OUT6_Mn6@78_d N_OUT5_Mn6@78_g N_VSS_Mn6@78_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@77 N_OUT6_Mn6@77_d N_OUT5_Mn6@77_g N_VSS_Mn6@77_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@76 N_OUT6_Mn6@76_d N_OUT5_Mn6@76_g N_VSS_Mn6@76_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@75 N_OUT6_Mn6@75_d N_OUT5_Mn6@75_g N_VSS_Mn6@75_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@74 N_OUT6_Mn6@74_d N_OUT5_Mn6@74_g N_VSS_Mn6@74_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@73 N_OUT6_Mn6@73_d N_OUT5_Mn6@73_g N_VSS_Mn6@73_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@72 N_OUT6_Mn6@72_d N_OUT5_Mn6@72_g N_VSS_Mn6@72_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@71 N_OUT6_Mn6@71_d N_OUT5_Mn6@71_g N_VSS_Mn6@71_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@70 N_OUT6_Mn6@70_d N_OUT5_Mn6@70_g N_VSS_Mn6@70_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@69 N_OUT6_Mn6@69_d N_OUT5_Mn6@69_g N_VSS_Mn6@69_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@68 N_OUT6_Mn6@68_d N_OUT5_Mn6@68_g N_VSS_Mn6@68_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@67 N_OUT6_Mn6@67_d N_OUT5_Mn6@67_g N_VSS_Mn6@67_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@66 N_OUT6_Mn6@66_d N_OUT5_Mn6@66_g N_VSS_Mn6@66_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@65 N_OUT6_Mn6@65_d N_OUT5_Mn6@65_g N_VSS_Mn6@65_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@64 N_OUT6_Mn6@64_d N_OUT5_Mn6@64_g N_VSS_Mn6@64_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@63 N_OUT6_Mn6@63_d N_OUT5_Mn6@63_g N_VSS_Mn6@63_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@62 N_OUT6_Mn6@62_d N_OUT5_Mn6@62_g N_VSS_Mn6@62_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@61 N_OUT6_Mn6@61_d N_OUT5_Mn6@61_g N_VSS_Mn6@61_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@60 N_OUT6_Mn6@60_d N_OUT5_Mn6@60_g N_VSS_Mn6@60_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@59 N_OUT6_Mn6@59_d N_OUT5_Mn6@59_g N_VSS_Mn6@59_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@58 N_OUT6_Mn6@58_d N_OUT5_Mn6@58_g N_VSS_Mn6@58_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@57 N_OUT6_Mn6@57_d N_OUT5_Mn6@57_g N_VSS_Mn6@57_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@56 N_OUT6_Mn6@56_d N_OUT5_Mn6@56_g N_VSS_Mn6@56_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@55 N_OUT6_Mn6@55_d N_OUT5_Mn6@55_g N_VSS_Mn6@55_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@54 N_OUT6_Mn6@54_d N_OUT5_Mn6@54_g N_VSS_Mn6@54_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@53 N_OUT6_Mn6@53_d N_OUT5_Mn6@53_g N_VSS_Mn6@53_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@52 N_OUT6_Mn6@52_d N_OUT5_Mn6@52_g N_VSS_Mn6@52_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@51 N_OUT6_Mn6@51_d N_OUT5_Mn6@51_g N_VSS_Mn6@51_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@50 N_OUT6_Mn6@50_d N_OUT5_Mn6@50_g N_VSS_Mn6@50_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@49 N_OUT6_Mn6@49_d N_OUT5_Mn6@49_g N_VSS_Mn6@49_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@48 N_OUT6_Mn6@48_d N_OUT5_Mn6@48_g N_VSS_Mn6@48_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@47 N_OUT6_Mn6@47_d N_OUT5_Mn6@47_g N_VSS_Mn6@47_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@46 N_OUT6_Mn6@46_d N_OUT5_Mn6@46_g N_VSS_Mn6@46_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@45 N_OUT6_Mn6@45_d N_OUT5_Mn6@45_g N_VSS_Mn6@45_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@44 N_OUT6_Mn6@44_d N_OUT5_Mn6@44_g N_VSS_Mn6@44_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@43 N_OUT6_Mn6@43_d N_OUT5_Mn6@43_g N_VSS_Mn6@43_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@42 N_OUT6_Mn6@42_d N_OUT5_Mn6@42_g N_VSS_Mn6@42_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@41 N_OUT6_Mn6@41_d N_OUT5_Mn6@41_g N_VSS_Mn6@41_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@40 N_OUT6_Mn6@40_d N_OUT5_Mn6@40_g N_VSS_Mn6@40_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@39 N_OUT6_Mn6@39_d N_OUT5_Mn6@39_g N_VSS_Mn6@39_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@38 N_OUT6_Mn6@38_d N_OUT5_Mn6@38_g N_VSS_Mn6@38_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@37 N_OUT6_Mn6@37_d N_OUT5_Mn6@37_g N_VSS_Mn6@37_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@36 N_OUT6_Mn6@36_d N_OUT5_Mn6@36_g N_VSS_Mn6@36_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@35 N_OUT6_Mn6@35_d N_OUT5_Mn6@35_g N_VSS_Mn6@35_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@34 N_OUT6_Mn6@34_d N_OUT5_Mn6@34_g N_VSS_Mn6@34_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@33 N_OUT6_Mn6@33_d N_OUT5_Mn6@33_g N_VSS_Mn6@33_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@32 N_OUT6_Mn6@32_d N_OUT5_Mn6@32_g N_VSS_Mn6@32_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@31 N_OUT6_Mn6@31_d N_OUT5_Mn6@31_g N_VSS_Mn6@31_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@30 N_OUT6_Mn6@30_d N_OUT5_Mn6@30_g N_VSS_Mn6@30_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@29 N_OUT6_Mn6@29_d N_OUT5_Mn6@29_g N_VSS_Mn6@29_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@28 N_OUT6_Mn6@28_d N_OUT5_Mn6@28_g N_VSS_Mn6@28_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@27 N_OUT6_Mn6@27_d N_OUT5_Mn6@27_g N_VSS_Mn6@27_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@26 N_OUT6_Mn6@26_d N_OUT5_Mn6@26_g N_VSS_Mn6@26_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@25 N_OUT6_Mn6@25_d N_OUT5_Mn6@25_g N_VSS_Mn6@25_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@24 N_OUT6_Mn6@24_d N_OUT5_Mn6@24_g N_VSS_Mn6@24_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@23 N_OUT6_Mn6@23_d N_OUT5_Mn6@23_g N_VSS_Mn6@23_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@22 N_OUT6_Mn6@22_d N_OUT5_Mn6@22_g N_VSS_Mn6@22_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@21 N_OUT6_Mn6@21_d N_OUT5_Mn6@21_g N_VSS_Mn6@21_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@20 N_OUT6_Mn6@20_d N_OUT5_Mn6@20_g N_VSS_Mn6@20_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@19 N_OUT6_Mn6@19_d N_OUT5_Mn6@19_g N_VSS_Mn6@19_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@18 N_OUT6_Mn6@18_d N_OUT5_Mn6@18_g N_VSS_Mn6@18_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@17 N_OUT6_Mn6@17_d N_OUT5_Mn6@17_g N_VSS_Mn6@17_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@16 N_OUT6_Mn6@16_d N_OUT5_Mn6@16_g N_VSS_Mn6@16_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@15 N_OUT6_Mn6@15_d N_OUT5_Mn6@15_g N_VSS_Mn6@15_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@14 N_OUT6_Mn6@14_d N_OUT5_Mn6@14_g N_VSS_Mn6@14_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@13 N_OUT6_Mn6@13_d N_OUT5_Mn6@13_g N_VSS_Mn6@13_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@12 N_OUT6_Mn6@12_d N_OUT5_Mn6@12_g N_VSS_Mn6@12_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@11 N_OUT6_Mn6@11_d N_OUT5_Mn6@11_g N_VSS_Mn6@11_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@10 N_OUT6_Mn6@10_d N_OUT5_Mn6@10_g N_VSS_Mn6@10_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@9 N_OUT6_Mn6@9_d N_OUT5_Mn6@9_g N_VSS_Mn6@9_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@8 N_OUT6_Mn6@8_d N_OUT5_Mn6@8_g N_VSS_Mn6@8_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@7 N_OUT6_Mn6@7_d N_OUT5_Mn6@7_g N_VSS_Mn6@7_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@6 N_OUT6_Mn6@6_d N_OUT5_Mn6@6_g N_VSS_Mn6@6_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@5 N_OUT6_Mn6@5_d N_OUT5_Mn6@5_g N_VSS_Mn6@5_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@4 N_OUT6_Mn6@4_d N_OUT5_Mn6@4_g N_VSS_Mn6@4_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@3 N_OUT6_Mn6@3_d N_OUT5_Mn6@3_g N_VSS_Mn6@3_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn6@2 N_OUT6_Mn6@2_d N_OUT5_Mn6@2_g N_VSS_Mn6@2_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=2.955e-13 AS=1.4125e-13 PD=1.682e-06 PS=5.65e-07
Mn7 N_OUT7_Mn7_d N_OUT6_Mn7_g N_VSS_Mn7_s N_VSS_Mn7@1159_b N_18 L=1.8e-07
+ W=5e-07 AD=1.325e-13 AS=2.995e-13 PD=5.3e-07 PS=1.698e-06
Mn7@1163 N_OUT7_Mn7@1163_d N_OUT6_Mn7@1163_g N_VSS_Mn7@1163_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1162 N_OUT7_Mn7@1162_d N_OUT6_Mn7@1162_g N_VSS_Mn7@1162_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1161 N_OUT7_Mn7@1161_d N_OUT6_Mn7@1161_g N_VSS_Mn7@1161_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1160 N_OUT7_Mn7@1160_d N_OUT6_Mn7@1160_g N_VSS_Mn7@1160_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.955e-13 AS=1.4125e-13 PD=1.682e-06 PS=5.65e-07
Mn8 N_OUT8_Mn8_d N_OUT7_Mn8_g N_VSS_Mn8_s N_VSS_Mn7@1159_b N_18 L=1.8e-07
+ W=5e-07 AD=1.325e-13 AS=2.995e-13 PD=5.3e-07 PS=1.698e-06
Mn8@3773 N_OUT8_Mn8@3773_d N_OUT7_Mn8@3773_g N_VSS_Mn8@3773_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3772 N_OUT8_Mn8@3772_d N_OUT7_Mn8@3772_g N_VSS_Mn8@3772_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3771 N_OUT8_Mn8@3771_d N_OUT7_Mn8@3771_g N_VSS_Mn8@3771_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4999 N_OUT9_Mn9@4999_d N_OUT8_Mn9@4999_g N_VSS_Mn9@4999_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4998 N_OUT9_Mn9@4998_d N_OUT8_Mn9@4998_g N_VSS_Mn9@4998_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4997 N_OUT9_Mn9@4997_d N_OUT8_Mn9@4997_g N_VSS_Mn9@4997_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4996 N_OUT9_Mn9@4996_d N_OUT8_Mn9@4996_g N_VSS_Mn9@4996_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=6.589e-13 PD=5.3e-07 PS=2.298e-06
Mn8@3770 N_OUT8_Mn8@3770_d N_OUT7_Mn8@3770_g N_VSS_Mn8@3770_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.955e-13 AS=1.4125e-13 PD=1.682e-06 PS=5.65e-07
Mp1 N_OUT1_Mp1_d N_OUT9_Mp1_g N_VDD_Mp1_s N_VDD_Mp1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.575e-13 AS=7.575e-13 PD=2.51e-06 PS=2.51e-06
Mp2 N_OUT2_Mp2_d N_OUT1_Mp2_g N_VDD_Mp2_s N_VDD_Mp2_b P_18 L=1.8e-07 W=1.5e-06
+ AD=3.9375e-13 AS=7.575e-13 PD=5.25e-07 PS=2.51e-06
Mp2@3 N_OUT2_Mp2@3_d N_OUT1_Mp2@3_g N_VDD_Mp2@3_s N_VDD_Mp2_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=3.9375e-13 PD=5.25e-07 PS=5.25e-07
Mp2@2 N_OUT2_Mp2@2_d N_OUT1_Mp2@2_g N_VDD_Mp2@2_s N_VDD_Mp2_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.575e-13 AS=3.9375e-13 PD=2.51e-06 PS=5.25e-07
Mp3 N_OUT3_Mp3_d N_OUT2_Mp3_g N_VDD_Mp3_s N_VDD_Mp3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=3.9375e-13 AS=7.575e-13 PD=5.25e-07 PS=2.51e-06
Mp3@11 N_OUT3_Mp3@11_d N_OUT2_Mp3@11_g N_VDD_Mp3@11_s N_VDD_Mp3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp3@10 N_OUT3_Mp3@10_d N_OUT2_Mp3@10_g N_VDD_Mp3@10_s N_VDD_Mp3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp3@9 N_OUT3_Mp3@9_d N_OUT2_Mp3@9_g N_VDD_Mp3@9_s N_VDD_Mp3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp3@8 N_OUT3_Mp3@8_d N_OUT2_Mp3@8_g N_VDD_Mp3@8_s N_VDD_Mp3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp3@7 N_OUT3_Mp3@7_d N_OUT2_Mp3@7_g N_VDD_Mp3@7_s N_VDD_Mp3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp3@6 N_OUT3_Mp3@6_d N_OUT2_Mp3@6_g N_VDD_Mp3@6_s N_VDD_Mp3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp3@5 N_OUT3_Mp3@5_d N_OUT2_Mp3@5_g N_VDD_Mp3@5_s N_VDD_Mp3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp3@4 N_OUT3_Mp3@4_d N_OUT2_Mp3@4_g N_VDD_Mp3@4_s N_VDD_Mp3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp3@3 N_OUT3_Mp3@3_d N_OUT2_Mp3@3_g N_VDD_Mp3@3_s N_VDD_Mp3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp3@2 N_OUT3_Mp3@2_d N_OUT2_Mp3@2_g N_VDD_Mp3@2_s N_VDD_Mp3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.575e-13 AS=4.275e-13 PD=2.51e-06 PS=5.7e-07
Mp4 N_OUT4_Mp4_d N_OUT3_Mp4_g N_VDD_Mp4_s N_VDD_Mp4_b P_18 L=1.8e-07 W=1.5e-06
+ AD=3.9375e-13 AS=7.575e-13 PD=5.25e-07 PS=2.51e-06
Mp4@34 N_OUT4_Mp4@34_d N_OUT3_Mp4@34_g N_VDD_Mp4@34_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@33 N_OUT4_Mp4@33_d N_OUT3_Mp4@33_g N_VDD_Mp4@33_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@32 N_OUT4_Mp4@32_d N_OUT3_Mp4@32_g N_VDD_Mp4@32_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@31 N_OUT4_Mp4@31_d N_OUT3_Mp4@31_g N_VDD_Mp4@31_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@30 N_OUT4_Mp4@30_d N_OUT3_Mp4@30_g N_VDD_Mp4@30_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@29 N_OUT4_Mp4@29_d N_OUT3_Mp4@29_g N_VDD_Mp4@29_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@28 N_OUT4_Mp4@28_d N_OUT3_Mp4@28_g N_VDD_Mp4@28_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@27 N_OUT4_Mp4@27_d N_OUT3_Mp4@27_g N_VDD_Mp4@27_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@26 N_OUT4_Mp4@26_d N_OUT3_Mp4@26_g N_VDD_Mp4@26_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@25 N_OUT4_Mp4@25_d N_OUT3_Mp4@25_g N_VDD_Mp4@25_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@24 N_OUT4_Mp4@24_d N_OUT3_Mp4@24_g N_VDD_Mp4@24_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@23 N_OUT4_Mp4@23_d N_OUT3_Mp4@23_g N_VDD_Mp4@23_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@22 N_OUT4_Mp4@22_d N_OUT3_Mp4@22_g N_VDD_Mp4@22_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@21 N_OUT4_Mp4@21_d N_OUT3_Mp4@21_g N_VDD_Mp4@21_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@20 N_OUT4_Mp4@20_d N_OUT3_Mp4@20_g N_VDD_Mp4@20_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@19 N_OUT4_Mp4@19_d N_OUT3_Mp4@19_g N_VDD_Mp4@19_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@18 N_OUT4_Mp4@18_d N_OUT3_Mp4@18_g N_VDD_Mp4@18_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@17 N_OUT4_Mp4@17_d N_OUT3_Mp4@17_g N_VDD_Mp4@17_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@16 N_OUT4_Mp4@16_d N_OUT3_Mp4@16_g N_VDD_Mp4@16_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@15 N_OUT4_Mp4@15_d N_OUT3_Mp4@15_g N_VDD_Mp4@15_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@14 N_OUT4_Mp4@14_d N_OUT3_Mp4@14_g N_VDD_Mp4@14_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@13 N_OUT4_Mp4@13_d N_OUT3_Mp4@13_g N_VDD_Mp4@13_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@12 N_OUT4_Mp4@12_d N_OUT3_Mp4@12_g N_VDD_Mp4@12_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@11 N_OUT4_Mp4@11_d N_OUT3_Mp4@11_g N_VDD_Mp4@11_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@10 N_OUT4_Mp4@10_d N_OUT3_Mp4@10_g N_VDD_Mp4@10_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@9 N_OUT4_Mp4@9_d N_OUT3_Mp4@9_g N_VDD_Mp4@9_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@8 N_OUT4_Mp4@8_d N_OUT3_Mp4@8_g N_VDD_Mp4@8_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@7 N_OUT4_Mp4@7_d N_OUT3_Mp4@7_g N_VDD_Mp4@7_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@6 N_OUT4_Mp4@6_d N_OUT3_Mp4@6_g N_VDD_Mp4@6_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@5 N_OUT4_Mp4@5_d N_OUT3_Mp4@5_g N_VDD_Mp4@5_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp4@4 N_OUT4_Mp4@4_d N_OUT3_Mp4@4_g N_VDD_Mp4@4_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=3.9375e-13 PD=5.25e-07 PS=5.25e-07
Mp4@3 N_OUT4_Mp4@3_d N_OUT3_Mp4@3_g N_VDD_Mp4@3_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=4.2e-13 AS=3.9375e-13 PD=5.6e-07 PS=5.25e-07
Mp4@2 N_OUT4_Mp4@2_d N_OUT3_Mp4@2_g N_VDD_Mp4@2_s N_VDD_Mp4_b P_18 L=1.8e-07
+ W=1.5e-06 AD=4.2e-13 AS=7.575e-13 PD=5.6e-07 PS=2.51e-06
Mp5 N_OUT5_Mp5_d N_OUT4_Mp5_g N_VDD_Mp5_s N_VDD_Mp5@105_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=7.575e-13 PD=5.25e-07 PS=2.51e-06
Mp5@111 N_OUT5_Mp5@111_d N_OUT4_Mp5@111_g N_VDD_Mp5@111_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@110 N_OUT5_Mp5@110_d N_OUT4_Mp5@110_g N_VDD_Mp5@110_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@109 N_OUT5_Mp5@109_d N_OUT4_Mp5@109_g N_VDD_Mp5@109_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@108 N_OUT5_Mp5@108_d N_OUT4_Mp5@108_g N_VDD_Mp5@108_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@107 N_OUT5_Mp5@107_d N_OUT4_Mp5@107_g N_VDD_Mp5@107_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@106 N_OUT5_Mp5@106_d N_OUT4_Mp5@106_g N_VDD_Mp5@106_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.575e-13 AS=4.275e-13 PD=2.51e-06 PS=5.7e-07
Mp6 N_OUT6_Mp6_d N_OUT5_Mp6_g N_VDD_Mp6_s N_VDD_Mp6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=3.9375e-13 AS=7.575e-13 PD=5.25e-07 PS=2.51e-06
Mp9 N_OUT9_Mp9_d N_OUT8_Mp9_g N_VDD_Mp9_s N_VDD_Mp9@4995_b P_18 L=1.8e-07
+ W=3.3e-06 AD=1.6665e-12 AS=9.405e-13 PD=4.31e-06 PS=5.7e-07
Mp6@359 N_OUT6_Mp6@359_d N_OUT5_Mp6@359_g N_VDD_Mp6@359_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@358 N_OUT6_Mp6@358_d N_OUT5_Mp6@358_g N_VDD_Mp6@358_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@357 N_OUT6_Mp6@357_d N_OUT5_Mp6@357_g N_VDD_Mp6@357_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@356 N_OUT6_Mp6@356_d N_OUT5_Mp6@356_g N_VDD_Mp6@356_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@355 N_OUT6_Mp6@355_d N_OUT5_Mp6@355_g N_VDD_Mp6@355_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@354 N_OUT6_Mp6@354_d N_OUT5_Mp6@354_g N_VDD_Mp6@354_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@353 N_OUT6_Mp6@353_d N_OUT5_Mp6@353_g N_VDD_Mp6@353_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@352 N_OUT6_Mp6@352_d N_OUT5_Mp6@352_g N_VDD_Mp6@352_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@351 N_OUT6_Mp6@351_d N_OUT5_Mp6@351_g N_VDD_Mp6@351_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@350 N_OUT6_Mp6@350_d N_OUT5_Mp6@350_g N_VDD_Mp6@350_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@349 N_OUT6_Mp6@349_d N_OUT5_Mp6@349_g N_VDD_Mp6@349_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@348 N_OUT6_Mp6@348_d N_OUT5_Mp6@348_g N_VDD_Mp6@348_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@347 N_OUT6_Mp6@347_d N_OUT5_Mp6@347_g N_VDD_Mp6@347_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@346 N_OUT6_Mp6@346_d N_OUT5_Mp6@346_g N_VDD_Mp6@346_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@345 N_OUT6_Mp6@345_d N_OUT5_Mp6@345_g N_VDD_Mp6@345_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@344 N_OUT6_Mp6@344_d N_OUT5_Mp6@344_g N_VDD_Mp6@344_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@343 N_OUT6_Mp6@343_d N_OUT5_Mp6@343_g N_VDD_Mp6@343_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@342 N_OUT6_Mp6@342_d N_OUT5_Mp6@342_g N_VDD_Mp6@342_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@341 N_OUT6_Mp6@341_d N_OUT5_Mp6@341_g N_VDD_Mp6@341_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@340 N_OUT6_Mp6@340_d N_OUT5_Mp6@340_g N_VDD_Mp6@340_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@339 N_OUT6_Mp6@339_d N_OUT5_Mp6@339_g N_VDD_Mp6@339_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@338 N_OUT6_Mp6@338_d N_OUT5_Mp6@338_g N_VDD_Mp6@338_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@337 N_OUT6_Mp6@337_d N_OUT5_Mp6@337_g N_VDD_Mp6@337_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@336 N_OUT6_Mp6@336_d N_OUT5_Mp6@336_g N_VDD_Mp6@336_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@335 N_OUT6_Mp6@335_d N_OUT5_Mp6@335_g N_VDD_Mp6@335_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@334 N_OUT6_Mp6@334_d N_OUT5_Mp6@334_g N_VDD_Mp6@334_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@333 N_OUT6_Mp6@333_d N_OUT5_Mp6@333_g N_VDD_Mp6@333_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@332 N_OUT6_Mp6@332_d N_OUT5_Mp6@332_g N_VDD_Mp6@332_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@331 N_OUT6_Mp6@331_d N_OUT5_Mp6@331_g N_VDD_Mp6@331_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@330 N_OUT6_Mp6@330_d N_OUT5_Mp6@330_g N_VDD_Mp6@330_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@329 N_OUT6_Mp6@329_d N_OUT5_Mp6@329_g N_VDD_Mp6@329_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@328 N_OUT6_Mp6@328_d N_OUT5_Mp6@328_g N_VDD_Mp6@328_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@327 N_OUT6_Mp6@327_d N_OUT5_Mp6@327_g N_VDD_Mp6@327_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@326 N_OUT6_Mp6@326_d N_OUT5_Mp6@326_g N_VDD_Mp6@326_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@325 N_OUT6_Mp6@325_d N_OUT5_Mp6@325_g N_VDD_Mp6@325_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@324 N_OUT6_Mp6@324_d N_OUT5_Mp6@324_g N_VDD_Mp6@324_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@323 N_OUT6_Mp6@323_d N_OUT5_Mp6@323_g N_VDD_Mp6@323_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@322 N_OUT6_Mp6@322_d N_OUT5_Mp6@322_g N_VDD_Mp6@322_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@321 N_OUT6_Mp6@321_d N_OUT5_Mp6@321_g N_VDD_Mp6@321_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@320 N_OUT6_Mp6@320_d N_OUT5_Mp6@320_g N_VDD_Mp6@320_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@319 N_OUT6_Mp6@319_d N_OUT5_Mp6@319_g N_VDD_Mp6@319_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@318 N_OUT6_Mp6@318_d N_OUT5_Mp6@318_g N_VDD_Mp6@318_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@317 N_OUT6_Mp6@317_d N_OUT5_Mp6@317_g N_VDD_Mp6@317_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@316 N_OUT6_Mp6@316_d N_OUT5_Mp6@316_g N_VDD_Mp6@316_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@315 N_OUT6_Mp6@315_d N_OUT5_Mp6@315_g N_VDD_Mp6@315_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@314 N_OUT6_Mp6@314_d N_OUT5_Mp6@314_g N_VDD_Mp6@314_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@313 N_OUT6_Mp6@313_d N_OUT5_Mp6@313_g N_VDD_Mp6@313_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@312 N_OUT6_Mp6@312_d N_OUT5_Mp6@312_g N_VDD_Mp6@312_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@311 N_OUT6_Mp6@311_d N_OUT5_Mp6@311_g N_VDD_Mp6@311_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@310 N_OUT6_Mp6@310_d N_OUT5_Mp6@310_g N_VDD_Mp6@310_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@309 N_OUT6_Mp6@309_d N_OUT5_Mp6@309_g N_VDD_Mp6@309_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@308 N_OUT6_Mp6@308_d N_OUT5_Mp6@308_g N_VDD_Mp6@308_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@307 N_OUT6_Mp6@307_d N_OUT5_Mp6@307_g N_VDD_Mp6@307_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@306 N_OUT6_Mp6@306_d N_OUT5_Mp6@306_g N_VDD_Mp6@306_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@305 N_OUT6_Mp6@305_d N_OUT5_Mp6@305_g N_VDD_Mp6@305_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@304 N_OUT6_Mp6@304_d N_OUT5_Mp6@304_g N_VDD_Mp6@304_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@303 N_OUT6_Mp6@303_d N_OUT5_Mp6@303_g N_VDD_Mp6@303_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@302 N_OUT6_Mp6@302_d N_OUT5_Mp6@302_g N_VDD_Mp6@302_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@301 N_OUT6_Mp6@301_d N_OUT5_Mp6@301_g N_VDD_Mp6@301_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@300 N_OUT6_Mp6@300_d N_OUT5_Mp6@300_g N_VDD_Mp6@300_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@299 N_OUT6_Mp6@299_d N_OUT5_Mp6@299_g N_VDD_Mp6@299_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@298 N_OUT6_Mp6@298_d N_OUT5_Mp6@298_g N_VDD_Mp6@298_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@297 N_OUT6_Mp6@297_d N_OUT5_Mp6@297_g N_VDD_Mp6@297_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@296 N_OUT6_Mp6@296_d N_OUT5_Mp6@296_g N_VDD_Mp6@296_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@295 N_OUT6_Mp6@295_d N_OUT5_Mp6@295_g N_VDD_Mp6@295_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@294 N_OUT6_Mp6@294_d N_OUT5_Mp6@294_g N_VDD_Mp6@294_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@293 N_OUT6_Mp6@293_d N_OUT5_Mp6@293_g N_VDD_Mp6@293_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@292 N_OUT6_Mp6@292_d N_OUT5_Mp6@292_g N_VDD_Mp6@292_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@291 N_OUT6_Mp6@291_d N_OUT5_Mp6@291_g N_VDD_Mp6@291_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@290 N_OUT6_Mp6@290_d N_OUT5_Mp6@290_g N_VDD_Mp6@290_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@289 N_OUT6_Mp6@289_d N_OUT5_Mp6@289_g N_VDD_Mp6@289_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@288 N_OUT6_Mp6@288_d N_OUT5_Mp6@288_g N_VDD_Mp6@288_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@287 N_OUT6_Mp6@287_d N_OUT5_Mp6@287_g N_VDD_Mp6@287_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@286 N_OUT6_Mp6@286_d N_OUT5_Mp6@286_g N_VDD_Mp6@286_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@285 N_OUT6_Mp6@285_d N_OUT5_Mp6@285_g N_VDD_Mp6@285_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@284 N_OUT6_Mp6@284_d N_OUT5_Mp6@284_g N_VDD_Mp6@284_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@283 N_OUT6_Mp6@283_d N_OUT5_Mp6@283_g N_VDD_Mp6@283_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@282 N_OUT6_Mp6@282_d N_OUT5_Mp6@282_g N_VDD_Mp6@282_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@281 N_OUT6_Mp6@281_d N_OUT5_Mp6@281_g N_VDD_Mp6@281_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@280 N_OUT6_Mp6@280_d N_OUT5_Mp6@280_g N_VDD_Mp6@280_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@279 N_OUT6_Mp6@279_d N_OUT5_Mp6@279_g N_VDD_Mp6@279_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@278 N_OUT6_Mp6@278_d N_OUT5_Mp6@278_g N_VDD_Mp6@278_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@277 N_OUT6_Mp6@277_d N_OUT5_Mp6@277_g N_VDD_Mp6@277_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@276 N_OUT6_Mp6@276_d N_OUT5_Mp6@276_g N_VDD_Mp6@276_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@275 N_OUT6_Mp6@275_d N_OUT5_Mp6@275_g N_VDD_Mp6@275_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@274 N_OUT6_Mp6@274_d N_OUT5_Mp6@274_g N_VDD_Mp6@274_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@273 N_OUT6_Mp6@273_d N_OUT5_Mp6@273_g N_VDD_Mp6@273_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@272 N_OUT6_Mp6@272_d N_OUT5_Mp6@272_g N_VDD_Mp6@272_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@271 N_OUT6_Mp6@271_d N_OUT5_Mp6@271_g N_VDD_Mp6@271_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@270 N_OUT6_Mp6@270_d N_OUT5_Mp6@270_g N_VDD_Mp6@270_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@269 N_OUT6_Mp6@269_d N_OUT5_Mp6@269_g N_VDD_Mp6@269_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@268 N_OUT6_Mp6@268_d N_OUT5_Mp6@268_g N_VDD_Mp6@268_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@267 N_OUT6_Mp6@267_d N_OUT5_Mp6@267_g N_VDD_Mp6@267_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@266 N_OUT6_Mp6@266_d N_OUT5_Mp6@266_g N_VDD_Mp6@266_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@265 N_OUT6_Mp6@265_d N_OUT5_Mp6@265_g N_VDD_Mp6@265_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@264 N_OUT6_Mp6@264_d N_OUT5_Mp6@264_g N_VDD_Mp6@264_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@263 N_OUT6_Mp6@263_d N_OUT5_Mp6@263_g N_VDD_Mp6@263_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@262 N_OUT6_Mp6@262_d N_OUT5_Mp6@262_g N_VDD_Mp6@262_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@261 N_OUT6_Mp6@261_d N_OUT5_Mp6@261_g N_VDD_Mp6@261_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@260 N_OUT6_Mp6@260_d N_OUT5_Mp6@260_g N_VDD_Mp6@260_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@259 N_OUT6_Mp6@259_d N_OUT5_Mp6@259_g N_VDD_Mp6@259_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@258 N_OUT6_Mp6@258_d N_OUT5_Mp6@258_g N_VDD_Mp6@258_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@257 N_OUT6_Mp6@257_d N_OUT5_Mp6@257_g N_VDD_Mp6@257_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@256 N_OUT6_Mp6@256_d N_OUT5_Mp6@256_g N_VDD_Mp6@256_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@255 N_OUT6_Mp6@255_d N_OUT5_Mp6@255_g N_VDD_Mp6@255_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@254 N_OUT6_Mp6@254_d N_OUT5_Mp6@254_g N_VDD_Mp6@254_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@253 N_OUT6_Mp6@253_d N_OUT5_Mp6@253_g N_VDD_Mp6@253_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@252 N_OUT6_Mp6@252_d N_OUT5_Mp6@252_g N_VDD_Mp6@252_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@251 N_OUT6_Mp6@251_d N_OUT5_Mp6@251_g N_VDD_Mp6@251_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@250 N_OUT6_Mp6@250_d N_OUT5_Mp6@250_g N_VDD_Mp6@250_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@249 N_OUT6_Mp6@249_d N_OUT5_Mp6@249_g N_VDD_Mp6@249_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@248 N_OUT6_Mp6@248_d N_OUT5_Mp6@248_g N_VDD_Mp6@248_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@247 N_OUT6_Mp6@247_d N_OUT5_Mp6@247_g N_VDD_Mp6@247_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@246 N_OUT6_Mp6@246_d N_OUT5_Mp6@246_g N_VDD_Mp6@246_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@245 N_OUT6_Mp6@245_d N_OUT5_Mp6@245_g N_VDD_Mp6@245_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@244 N_OUT6_Mp6@244_d N_OUT5_Mp6@244_g N_VDD_Mp6@244_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@243 N_OUT6_Mp6@243_d N_OUT5_Mp6@243_g N_VDD_Mp6@243_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@242 N_OUT6_Mp6@242_d N_OUT5_Mp6@242_g N_VDD_Mp6@242_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@241 N_OUT6_Mp6@241_d N_OUT5_Mp6@241_g N_VDD_Mp6@241_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@240 N_OUT6_Mp6@240_d N_OUT5_Mp6@240_g N_VDD_Mp6@240_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@239 N_OUT6_Mp6@239_d N_OUT5_Mp6@239_g N_VDD_Mp6@239_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@238 N_OUT6_Mp6@238_d N_OUT5_Mp6@238_g N_VDD_Mp6@238_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@237 N_OUT6_Mp6@237_d N_OUT5_Mp6@237_g N_VDD_Mp6@237_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@236 N_OUT6_Mp6@236_d N_OUT5_Mp6@236_g N_VDD_Mp6@236_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@235 N_OUT6_Mp6@235_d N_OUT5_Mp6@235_g N_VDD_Mp6@235_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@234 N_OUT6_Mp6@234_d N_OUT5_Mp6@234_g N_VDD_Mp6@234_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@233 N_OUT6_Mp6@233_d N_OUT5_Mp6@233_g N_VDD_Mp6@233_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@232 N_OUT6_Mp6@232_d N_OUT5_Mp6@232_g N_VDD_Mp6@232_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@231 N_OUT6_Mp6@231_d N_OUT5_Mp6@231_g N_VDD_Mp6@231_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@230 N_OUT6_Mp6@230_d N_OUT5_Mp6@230_g N_VDD_Mp6@230_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@229 N_OUT6_Mp6@229_d N_OUT5_Mp6@229_g N_VDD_Mp6@229_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@228 N_OUT6_Mp6@228_d N_OUT5_Mp6@228_g N_VDD_Mp6@228_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@227 N_OUT6_Mp6@227_d N_OUT5_Mp6@227_g N_VDD_Mp6@227_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@226 N_OUT6_Mp6@226_d N_OUT5_Mp6@226_g N_VDD_Mp6@226_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@225 N_OUT6_Mp6@225_d N_OUT5_Mp6@225_g N_VDD_Mp6@225_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@224 N_OUT6_Mp6@224_d N_OUT5_Mp6@224_g N_VDD_Mp6@224_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@223 N_OUT6_Mp6@223_d N_OUT5_Mp6@223_g N_VDD_Mp6@223_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@222 N_OUT6_Mp6@222_d N_OUT5_Mp6@222_g N_VDD_Mp6@222_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@221 N_OUT6_Mp6@221_d N_OUT5_Mp6@221_g N_VDD_Mp6@221_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@220 N_OUT6_Mp6@220_d N_OUT5_Mp6@220_g N_VDD_Mp6@220_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@219 N_OUT6_Mp6@219_d N_OUT5_Mp6@219_g N_VDD_Mp6@219_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@218 N_OUT6_Mp6@218_d N_OUT5_Mp6@218_g N_VDD_Mp6@218_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@217 N_OUT6_Mp6@217_d N_OUT5_Mp6@217_g N_VDD_Mp6@217_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@216 N_OUT6_Mp6@216_d N_OUT5_Mp6@216_g N_VDD_Mp6@216_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@215 N_OUT6_Mp6@215_d N_OUT5_Mp6@215_g N_VDD_Mp6@215_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@214 N_OUT6_Mp6@214_d N_OUT5_Mp6@214_g N_VDD_Mp6@214_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@213 N_OUT6_Mp6@213_d N_OUT5_Mp6@213_g N_VDD_Mp6@213_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@212 N_OUT6_Mp6@212_d N_OUT5_Mp6@212_g N_VDD_Mp6@212_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@211 N_OUT6_Mp6@211_d N_OUT5_Mp6@211_g N_VDD_Mp6@211_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@210 N_OUT6_Mp6@210_d N_OUT5_Mp6@210_g N_VDD_Mp6@210_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@209 N_OUT6_Mp6@209_d N_OUT5_Mp6@209_g N_VDD_Mp6@209_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@208 N_OUT6_Mp6@208_d N_OUT5_Mp6@208_g N_VDD_Mp6@208_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@207 N_OUT6_Mp6@207_d N_OUT5_Mp6@207_g N_VDD_Mp6@207_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@206 N_OUT6_Mp6@206_d N_OUT5_Mp6@206_g N_VDD_Mp6@206_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@205 N_OUT6_Mp6@205_d N_OUT5_Mp6@205_g N_VDD_Mp6@205_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@204 N_OUT6_Mp6@204_d N_OUT5_Mp6@204_g N_VDD_Mp6@204_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@203 N_OUT6_Mp6@203_d N_OUT5_Mp6@203_g N_VDD_Mp6@203_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@202 N_OUT6_Mp6@202_d N_OUT5_Mp6@202_g N_VDD_Mp6@202_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@201 N_OUT6_Mp6@201_d N_OUT5_Mp6@201_g N_VDD_Mp6@201_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@200 N_OUT6_Mp6@200_d N_OUT5_Mp6@200_g N_VDD_Mp6@200_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@199 N_OUT6_Mp6@199_d N_OUT5_Mp6@199_g N_VDD_Mp6@199_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@198 N_OUT6_Mp6@198_d N_OUT5_Mp6@198_g N_VDD_Mp6@198_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@197 N_OUT6_Mp6@197_d N_OUT5_Mp6@197_g N_VDD_Mp6@197_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@196 N_OUT6_Mp6@196_d N_OUT5_Mp6@196_g N_VDD_Mp6@196_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@195 N_OUT6_Mp6@195_d N_OUT5_Mp6@195_g N_VDD_Mp6@195_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@194 N_OUT6_Mp6@194_d N_OUT5_Mp6@194_g N_VDD_Mp6@194_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@193 N_OUT6_Mp6@193_d N_OUT5_Mp6@193_g N_VDD_Mp6@193_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@192 N_OUT6_Mp6@192_d N_OUT5_Mp6@192_g N_VDD_Mp6@192_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@191 N_OUT6_Mp6@191_d N_OUT5_Mp6@191_g N_VDD_Mp6@191_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@190 N_OUT6_Mp6@190_d N_OUT5_Mp6@190_g N_VDD_Mp6@190_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@189 N_OUT6_Mp6@189_d N_OUT5_Mp6@189_g N_VDD_Mp6@189_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@188 N_OUT6_Mp6@188_d N_OUT5_Mp6@188_g N_VDD_Mp6@188_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@187 N_OUT6_Mp6@187_d N_OUT5_Mp6@187_g N_VDD_Mp6@187_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@186 N_OUT6_Mp6@186_d N_OUT5_Mp6@186_g N_VDD_Mp6@186_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@185 N_OUT6_Mp6@185_d N_OUT5_Mp6@185_g N_VDD_Mp6@185_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@184 N_OUT6_Mp6@184_d N_OUT5_Mp6@184_g N_VDD_Mp6@184_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@183 N_OUT6_Mp6@183_d N_OUT5_Mp6@183_g N_VDD_Mp6@183_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@182 N_OUT6_Mp6@182_d N_OUT5_Mp6@182_g N_VDD_Mp6@182_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@181 N_OUT6_Mp6@181_d N_OUT5_Mp6@181_g N_VDD_Mp6@181_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@180 N_OUT6_Mp6@180_d N_OUT5_Mp6@180_g N_VDD_Mp6@180_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@179 N_OUT6_Mp6@179_d N_OUT5_Mp6@179_g N_VDD_Mp6@179_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@178 N_OUT6_Mp6@178_d N_OUT5_Mp6@178_g N_VDD_Mp6@178_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@177 N_OUT6_Mp6@177_d N_OUT5_Mp6@177_g N_VDD_Mp6@177_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@176 N_OUT6_Mp6@176_d N_OUT5_Mp6@176_g N_VDD_Mp6@176_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@175 N_OUT6_Mp6@175_d N_OUT5_Mp6@175_g N_VDD_Mp6@175_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@174 N_OUT6_Mp6@174_d N_OUT5_Mp6@174_g N_VDD_Mp6@174_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@173 N_OUT6_Mp6@173_d N_OUT5_Mp6@173_g N_VDD_Mp6@173_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@172 N_OUT6_Mp6@172_d N_OUT5_Mp6@172_g N_VDD_Mp6@172_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@171 N_OUT6_Mp6@171_d N_OUT5_Mp6@171_g N_VDD_Mp6@171_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@170 N_OUT6_Mp6@170_d N_OUT5_Mp6@170_g N_VDD_Mp6@170_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@169 N_OUT6_Mp6@169_d N_OUT5_Mp6@169_g N_VDD_Mp6@169_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@168 N_OUT6_Mp6@168_d N_OUT5_Mp6@168_g N_VDD_Mp6@168_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@167 N_OUT6_Mp6@167_d N_OUT5_Mp6@167_g N_VDD_Mp6@167_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@166 N_OUT6_Mp6@166_d N_OUT5_Mp6@166_g N_VDD_Mp6@166_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@165 N_OUT6_Mp6@165_d N_OUT5_Mp6@165_g N_VDD_Mp6@165_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@164 N_OUT6_Mp6@164_d N_OUT5_Mp6@164_g N_VDD_Mp6@164_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@163 N_OUT6_Mp6@163_d N_OUT5_Mp6@163_g N_VDD_Mp6@163_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@162 N_OUT6_Mp6@162_d N_OUT5_Mp6@162_g N_VDD_Mp6@162_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@161 N_OUT6_Mp6@161_d N_OUT5_Mp6@161_g N_VDD_Mp6@161_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@160 N_OUT6_Mp6@160_d N_OUT5_Mp6@160_g N_VDD_Mp6@160_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@159 N_OUT6_Mp6@159_d N_OUT5_Mp6@159_g N_VDD_Mp6@159_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@158 N_OUT6_Mp6@158_d N_OUT5_Mp6@158_g N_VDD_Mp6@158_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@157 N_OUT6_Mp6@157_d N_OUT5_Mp6@157_g N_VDD_Mp6@157_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@156 N_OUT6_Mp6@156_d N_OUT5_Mp6@156_g N_VDD_Mp6@156_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@155 N_OUT6_Mp6@155_d N_OUT5_Mp6@155_g N_VDD_Mp6@155_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@154 N_OUT6_Mp6@154_d N_OUT5_Mp6@154_g N_VDD_Mp6@154_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@153 N_OUT6_Mp6@153_d N_OUT5_Mp6@153_g N_VDD_Mp6@153_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@152 N_OUT6_Mp6@152_d N_OUT5_Mp6@152_g N_VDD_Mp6@152_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@151 N_OUT6_Mp6@151_d N_OUT5_Mp6@151_g N_VDD_Mp6@151_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@150 N_OUT6_Mp6@150_d N_OUT5_Mp6@150_g N_VDD_Mp6@150_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@149 N_OUT6_Mp6@149_d N_OUT5_Mp6@149_g N_VDD_Mp6@149_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@148 N_OUT6_Mp6@148_d N_OUT5_Mp6@148_g N_VDD_Mp6@148_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@147 N_OUT6_Mp6@147_d N_OUT5_Mp6@147_g N_VDD_Mp6@147_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@146 N_OUT6_Mp6@146_d N_OUT5_Mp6@146_g N_VDD_Mp6@146_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@145 N_OUT6_Mp6@145_d N_OUT5_Mp6@145_g N_VDD_Mp6@145_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@144 N_OUT6_Mp6@144_d N_OUT5_Mp6@144_g N_VDD_Mp6@144_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@143 N_OUT6_Mp6@143_d N_OUT5_Mp6@143_g N_VDD_Mp6@143_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@142 N_OUT6_Mp6@142_d N_OUT5_Mp6@142_g N_VDD_Mp6@142_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@141 N_OUT6_Mp6@141_d N_OUT5_Mp6@141_g N_VDD_Mp6@141_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@140 N_OUT6_Mp6@140_d N_OUT5_Mp6@140_g N_VDD_Mp6@140_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@139 N_OUT6_Mp6@139_d N_OUT5_Mp6@139_g N_VDD_Mp6@139_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@138 N_OUT6_Mp6@138_d N_OUT5_Mp6@138_g N_VDD_Mp6@138_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@137 N_OUT6_Mp6@137_d N_OUT5_Mp6@137_g N_VDD_Mp6@137_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@136 N_OUT6_Mp6@136_d N_OUT5_Mp6@136_g N_VDD_Mp6@136_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@135 N_OUT6_Mp6@135_d N_OUT5_Mp6@135_g N_VDD_Mp6@135_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@134 N_OUT6_Mp6@134_d N_OUT5_Mp6@134_g N_VDD_Mp6@134_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@133 N_OUT6_Mp6@133_d N_OUT5_Mp6@133_g N_VDD_Mp6@133_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@132 N_OUT6_Mp6@132_d N_OUT5_Mp6@132_g N_VDD_Mp6@132_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@131 N_OUT6_Mp6@131_d N_OUT5_Mp6@131_g N_VDD_Mp6@131_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@130 N_OUT6_Mp6@130_d N_OUT5_Mp6@130_g N_VDD_Mp6@130_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@129 N_OUT6_Mp6@129_d N_OUT5_Mp6@129_g N_VDD_Mp6@129_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@128 N_OUT6_Mp6@128_d N_OUT5_Mp6@128_g N_VDD_Mp6@128_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@127 N_OUT6_Mp6@127_d N_OUT5_Mp6@127_g N_VDD_Mp6@127_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@126 N_OUT6_Mp6@126_d N_OUT5_Mp6@126_g N_VDD_Mp6@126_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@125 N_OUT6_Mp6@125_d N_OUT5_Mp6@125_g N_VDD_Mp6@125_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@124 N_OUT6_Mp6@124_d N_OUT5_Mp6@124_g N_VDD_Mp6@124_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@123 N_OUT6_Mp6@123_d N_OUT5_Mp6@123_g N_VDD_Mp6@123_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@122 N_OUT6_Mp6@122_d N_OUT5_Mp6@122_g N_VDD_Mp6@122_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@121 N_OUT6_Mp6@121_d N_OUT5_Mp6@121_g N_VDD_Mp6@121_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@120 N_OUT6_Mp6@120_d N_OUT5_Mp6@120_g N_VDD_Mp6@120_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@119 N_OUT6_Mp6@119_d N_OUT5_Mp6@119_g N_VDD_Mp6@119_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@118 N_OUT6_Mp6@118_d N_OUT5_Mp6@118_g N_VDD_Mp6@118_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@117 N_OUT6_Mp6@117_d N_OUT5_Mp6@117_g N_VDD_Mp6@117_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@116 N_OUT6_Mp6@116_d N_OUT5_Mp6@116_g N_VDD_Mp6@116_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@115 N_OUT6_Mp6@115_d N_OUT5_Mp6@115_g N_VDD_Mp6@115_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@114 N_OUT6_Mp6@114_d N_OUT5_Mp6@114_g N_VDD_Mp6@114_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@113 N_OUT6_Mp6@113_d N_OUT5_Mp6@113_g N_VDD_Mp6@113_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@112 N_OUT6_Mp6@112_d N_OUT5_Mp6@112_g N_VDD_Mp6@112_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@111 N_OUT6_Mp6@111_d N_OUT5_Mp6@111_g N_VDD_Mp6@111_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@110 N_OUT6_Mp6@110_d N_OUT5_Mp6@110_g N_VDD_Mp6@110_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@109 N_OUT6_Mp6@109_d N_OUT5_Mp6@109_g N_VDD_Mp6@109_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@108 N_OUT6_Mp6@108_d N_OUT5_Mp6@108_g N_VDD_Mp6@108_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@107 N_OUT6_Mp6@107_d N_OUT5_Mp6@107_g N_VDD_Mp6@107_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@106 N_OUT6_Mp6@106_d N_OUT5_Mp6@106_g N_VDD_Mp6@106_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@105 N_OUT6_Mp6@105_d N_OUT5_Mp6@105_g N_VDD_Mp6@105_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@104 N_OUT6_Mp6@104_d N_OUT5_Mp6@104_g N_VDD_Mp6@104_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@103 N_OUT6_Mp6@103_d N_OUT5_Mp6@103_g N_VDD_Mp6@103_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@102 N_OUT6_Mp6@102_d N_OUT5_Mp6@102_g N_VDD_Mp6@102_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@101 N_OUT6_Mp6@101_d N_OUT5_Mp6@101_g N_VDD_Mp6@101_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@100 N_OUT6_Mp6@100_d N_OUT5_Mp6@100_g N_VDD_Mp6@100_s N_VDD_Mp6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@99 N_OUT6_Mp6@99_d N_OUT5_Mp6@99_g N_VDD_Mp6@99_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@98 N_OUT6_Mp6@98_d N_OUT5_Mp6@98_g N_VDD_Mp6@98_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@97 N_OUT6_Mp6@97_d N_OUT5_Mp6@97_g N_VDD_Mp6@97_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@96 N_OUT6_Mp6@96_d N_OUT5_Mp6@96_g N_VDD_Mp6@96_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@95 N_OUT6_Mp6@95_d N_OUT5_Mp6@95_g N_VDD_Mp6@95_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@94 N_OUT6_Mp6@94_d N_OUT5_Mp6@94_g N_VDD_Mp6@94_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@93 N_OUT6_Mp6@93_d N_OUT5_Mp6@93_g N_VDD_Mp6@93_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@92 N_OUT6_Mp6@92_d N_OUT5_Mp6@92_g N_VDD_Mp6@92_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@91 N_OUT6_Mp6@91_d N_OUT5_Mp6@91_g N_VDD_Mp6@91_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@90 N_OUT6_Mp6@90_d N_OUT5_Mp6@90_g N_VDD_Mp6@90_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@89 N_OUT6_Mp6@89_d N_OUT5_Mp6@89_g N_VDD_Mp6@89_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@88 N_OUT6_Mp6@88_d N_OUT5_Mp6@88_g N_VDD_Mp6@88_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@87 N_OUT6_Mp6@87_d N_OUT5_Mp6@87_g N_VDD_Mp6@87_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@86 N_OUT6_Mp6@86_d N_OUT5_Mp6@86_g N_VDD_Mp6@86_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@85 N_OUT6_Mp6@85_d N_OUT5_Mp6@85_g N_VDD_Mp6@85_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@84 N_OUT6_Mp6@84_d N_OUT5_Mp6@84_g N_VDD_Mp6@84_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@83 N_OUT6_Mp6@83_d N_OUT5_Mp6@83_g N_VDD_Mp6@83_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@82 N_OUT6_Mp6@82_d N_OUT5_Mp6@82_g N_VDD_Mp6@82_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@81 N_OUT6_Mp6@81_d N_OUT5_Mp6@81_g N_VDD_Mp6@81_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@80 N_OUT6_Mp6@80_d N_OUT5_Mp6@80_g N_VDD_Mp6@80_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@79 N_OUT6_Mp6@79_d N_OUT5_Mp6@79_g N_VDD_Mp6@79_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@78 N_OUT6_Mp6@78_d N_OUT5_Mp6@78_g N_VDD_Mp6@78_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@77 N_OUT6_Mp6@77_d N_OUT5_Mp6@77_g N_VDD_Mp6@77_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@76 N_OUT6_Mp6@76_d N_OUT5_Mp6@76_g N_VDD_Mp6@76_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@75 N_OUT6_Mp6@75_d N_OUT5_Mp6@75_g N_VDD_Mp6@75_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@74 N_OUT6_Mp6@74_d N_OUT5_Mp6@74_g N_VDD_Mp6@74_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@73 N_OUT6_Mp6@73_d N_OUT5_Mp6@73_g N_VDD_Mp6@73_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@72 N_OUT6_Mp6@72_d N_OUT5_Mp6@72_g N_VDD_Mp6@72_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@71 N_OUT6_Mp6@71_d N_OUT5_Mp6@71_g N_VDD_Mp6@71_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@70 N_OUT6_Mp6@70_d N_OUT5_Mp6@70_g N_VDD_Mp6@70_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@69 N_OUT6_Mp6@69_d N_OUT5_Mp6@69_g N_VDD_Mp6@69_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@68 N_OUT6_Mp6@68_d N_OUT5_Mp6@68_g N_VDD_Mp6@68_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@67 N_OUT6_Mp6@67_d N_OUT5_Mp6@67_g N_VDD_Mp6@67_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@66 N_OUT6_Mp6@66_d N_OUT5_Mp6@66_g N_VDD_Mp6@66_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@65 N_OUT6_Mp6@65_d N_OUT5_Mp6@65_g N_VDD_Mp6@65_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@64 N_OUT6_Mp6@64_d N_OUT5_Mp6@64_g N_VDD_Mp6@64_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@63 N_OUT6_Mp6@63_d N_OUT5_Mp6@63_g N_VDD_Mp6@63_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@62 N_OUT6_Mp6@62_d N_OUT5_Mp6@62_g N_VDD_Mp6@62_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@61 N_OUT6_Mp6@61_d N_OUT5_Mp6@61_g N_VDD_Mp6@61_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@60 N_OUT6_Mp6@60_d N_OUT5_Mp6@60_g N_VDD_Mp6@60_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@59 N_OUT6_Mp6@59_d N_OUT5_Mp6@59_g N_VDD_Mp6@59_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@58 N_OUT6_Mp6@58_d N_OUT5_Mp6@58_g N_VDD_Mp6@58_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@57 N_OUT6_Mp6@57_d N_OUT5_Mp6@57_g N_VDD_Mp6@57_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@56 N_OUT6_Mp6@56_d N_OUT5_Mp6@56_g N_VDD_Mp6@56_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@55 N_OUT6_Mp6@55_d N_OUT5_Mp6@55_g N_VDD_Mp6@55_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@54 N_OUT6_Mp6@54_d N_OUT5_Mp6@54_g N_VDD_Mp6@54_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@53 N_OUT6_Mp6@53_d N_OUT5_Mp6@53_g N_VDD_Mp6@53_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@52 N_OUT6_Mp6@52_d N_OUT5_Mp6@52_g N_VDD_Mp6@52_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@51 N_OUT6_Mp6@51_d N_OUT5_Mp6@51_g N_VDD_Mp6@51_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@50 N_OUT6_Mp6@50_d N_OUT5_Mp6@50_g N_VDD_Mp6@50_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@49 N_OUT6_Mp6@49_d N_OUT5_Mp6@49_g N_VDD_Mp6@49_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@48 N_OUT6_Mp6@48_d N_OUT5_Mp6@48_g N_VDD_Mp6@48_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@47 N_OUT6_Mp6@47_d N_OUT5_Mp6@47_g N_VDD_Mp6@47_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@46 N_OUT6_Mp6@46_d N_OUT5_Mp6@46_g N_VDD_Mp6@46_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@45 N_OUT6_Mp6@45_d N_OUT5_Mp6@45_g N_VDD_Mp6@45_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@44 N_OUT6_Mp6@44_d N_OUT5_Mp6@44_g N_VDD_Mp6@44_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@43 N_OUT6_Mp6@43_d N_OUT5_Mp6@43_g N_VDD_Mp6@43_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@42 N_OUT6_Mp6@42_d N_OUT5_Mp6@42_g N_VDD_Mp6@42_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@41 N_OUT6_Mp6@41_d N_OUT5_Mp6@41_g N_VDD_Mp6@41_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@40 N_OUT6_Mp6@40_d N_OUT5_Mp6@40_g N_VDD_Mp6@40_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@39 N_OUT6_Mp6@39_d N_OUT5_Mp6@39_g N_VDD_Mp6@39_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@38 N_OUT6_Mp6@38_d N_OUT5_Mp6@38_g N_VDD_Mp6@38_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@37 N_OUT6_Mp6@37_d N_OUT5_Mp6@37_g N_VDD_Mp6@37_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@36 N_OUT6_Mp6@36_d N_OUT5_Mp6@36_g N_VDD_Mp6@36_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@35 N_OUT6_Mp6@35_d N_OUT5_Mp6@35_g N_VDD_Mp6@35_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@34 N_OUT6_Mp6@34_d N_OUT5_Mp6@34_g N_VDD_Mp6@34_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@33 N_OUT6_Mp6@33_d N_OUT5_Mp6@33_g N_VDD_Mp6@33_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@32 N_OUT6_Mp6@32_d N_OUT5_Mp6@32_g N_VDD_Mp6@32_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@31 N_OUT6_Mp6@31_d N_OUT5_Mp6@31_g N_VDD_Mp6@31_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@30 N_OUT6_Mp6@30_d N_OUT5_Mp6@30_g N_VDD_Mp6@30_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@29 N_OUT6_Mp6@29_d N_OUT5_Mp6@29_g N_VDD_Mp6@29_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@28 N_OUT6_Mp6@28_d N_OUT5_Mp6@28_g N_VDD_Mp6@28_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@27 N_OUT6_Mp6@27_d N_OUT5_Mp6@27_g N_VDD_Mp6@27_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@26 N_OUT6_Mp6@26_d N_OUT5_Mp6@26_g N_VDD_Mp6@26_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@25 N_OUT6_Mp6@25_d N_OUT5_Mp6@25_g N_VDD_Mp6@25_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@24 N_OUT6_Mp6@24_d N_OUT5_Mp6@24_g N_VDD_Mp6@24_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@23 N_OUT6_Mp6@23_d N_OUT5_Mp6@23_g N_VDD_Mp6@23_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@22 N_OUT6_Mp6@22_d N_OUT5_Mp6@22_g N_VDD_Mp6@22_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@21 N_OUT6_Mp6@21_d N_OUT5_Mp6@21_g N_VDD_Mp6@21_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@20 N_OUT6_Mp6@20_d N_OUT5_Mp6@20_g N_VDD_Mp6@20_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@19 N_OUT6_Mp6@19_d N_OUT5_Mp6@19_g N_VDD_Mp6@19_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@18 N_OUT6_Mp6@18_d N_OUT5_Mp6@18_g N_VDD_Mp6@18_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@17 N_OUT6_Mp6@17_d N_OUT5_Mp6@17_g N_VDD_Mp6@17_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@16 N_OUT6_Mp6@16_d N_OUT5_Mp6@16_g N_VDD_Mp6@16_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@15 N_OUT6_Mp6@15_d N_OUT5_Mp6@15_g N_VDD_Mp6@15_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@14 N_OUT6_Mp6@14_d N_OUT5_Mp6@14_g N_VDD_Mp6@14_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@13 N_OUT6_Mp6@13_d N_OUT5_Mp6@13_g N_VDD_Mp6@13_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@12 N_OUT6_Mp6@12_d N_OUT5_Mp6@12_g N_VDD_Mp6@12_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@11 N_OUT6_Mp6@11_d N_OUT5_Mp6@11_g N_VDD_Mp6@11_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@10 N_OUT6_Mp6@10_d N_OUT5_Mp6@10_g N_VDD_Mp6@10_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@9 N_OUT6_Mp6@9_d N_OUT5_Mp6@9_g N_VDD_Mp6@9_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@8 N_OUT6_Mp6@8_d N_OUT5_Mp6@8_g N_VDD_Mp6@8_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@7 N_OUT6_Mp6@7_d N_OUT5_Mp6@7_g N_VDD_Mp6@7_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@6 N_OUT6_Mp6@6_d N_OUT5_Mp6@6_g N_VDD_Mp6@6_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@5 N_OUT6_Mp6@5_d N_OUT5_Mp6@5_g N_VDD_Mp6@5_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@4 N_OUT6_Mp6@4_d N_OUT5_Mp6@4_g N_VDD_Mp6@4_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@3 N_OUT6_Mp6@3_d N_OUT5_Mp6@3_g N_VDD_Mp6@3_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp6@2 N_OUT6_Mp6@2_d N_OUT5_Mp6@2_g N_VDD_Mp6@2_s N_VDD_Mp6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.95e-13 AS=4.275e-13 PD=2.56e-06 PS=5.7e-07
Mp7 N_OUT7_Mp7_d N_OUT6_Mp7_g N_VDD_Mp7_s N_VDD_Mp7@1159_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=7.575e-13 PD=5.25e-07 PS=2.51e-06
Mp7@1163 N_OUT7_Mp7@1163_d N_OUT6_Mp7@1163_g N_VDD_Mp7@1163_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1162 N_OUT7_Mp7@1162_d N_OUT6_Mp7@1162_g N_VDD_Mp7@1162_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1161 N_OUT7_Mp7@1161_d N_OUT6_Mp7@1161_g N_VDD_Mp7@1161_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1160 N_OUT7_Mp7@1160_d N_OUT6_Mp7@1160_g N_VDD_Mp7@1160_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.575e-13 AS=4.275e-13 PD=2.51e-06 PS=5.7e-07
Mp8 N_OUT8_Mp8_d N_OUT7_Mp8_g N_VDD_Mp8_s N_VDD_Mp8@3769_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=7.575e-13 PD=5.25e-07 PS=2.51e-06
Mp8@3773 N_OUT8_Mp8@3773_d N_OUT7_Mp8@3773_g N_VDD_Mp8@3773_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3772 N_OUT8_Mp8@3772_d N_OUT7_Mp8@3772_g N_VDD_Mp8@3772_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3771 N_OUT8_Mp8@3771_d N_OUT7_Mp8@3771_g N_VDD_Mp8@3771_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4999 N_OUT9_Mp9@4999_d N_OUT8_Mp9@4999_g N_VDD_Mp9@4999_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4998 N_OUT9_Mp9@4998_d N_OUT8_Mp9@4998_g N_VDD_Mp9@4998_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4997 N_OUT9_Mp9@4997_d N_OUT8_Mp9@4997_g N_VDD_Mp9@4997_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4996 N_OUT9_Mp9@4996_d N_OUT8_Mp9@4996_g N_VDD_Mp9@4996_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=1.6665e-12 PD=5.25e-07 PS=4.31e-06
Mp8@3770 N_OUT8_Mp8@3770_d N_OUT7_Mp8@3770_g N_VDD_Mp8@3770_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.575e-13 AS=4.275e-13 PD=2.51e-06 PS=5.7e-07
Mn7@1159 N_OUT7_Mn7@1159_d N_OUT6_Mn7@1159_g N_VSS_Mn7@1159_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1158 N_OUT7_Mn7@1158_d N_OUT6_Mn7@1158_g N_VSS_Mn7@1158_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1159 N_OUT7_Mp7@1159_d N_OUT6_Mp7@1159_g N_VDD_Mp7@1159_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1158 N_OUT7_Mp7@1158_d N_OUT6_Mp7@1158_g N_VDD_Mp7@1158_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1157 N_OUT7_Mn7@1157_d N_OUT6_Mn7@1157_g N_VSS_Mn7@1157_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1156 N_OUT7_Mn7@1156_d N_OUT6_Mn7@1156_g N_VSS_Mn7@1156_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1157 N_OUT7_Mp7@1157_d N_OUT6_Mp7@1157_g N_VDD_Mp7@1157_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1156 N_OUT7_Mp7@1156_d N_OUT6_Mp7@1156_g N_VDD_Mp7@1156_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1155 N_OUT7_Mn7@1155_d N_OUT6_Mn7@1155_g N_VSS_Mn7@1155_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1154 N_OUT7_Mn7@1154_d N_OUT6_Mn7@1154_g N_VSS_Mn7@1154_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1155 N_OUT7_Mp7@1155_d N_OUT6_Mp7@1155_g N_VDD_Mp7@1155_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1154 N_OUT7_Mp7@1154_d N_OUT6_Mp7@1154_g N_VDD_Mp7@1154_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@105 N_OUT5_Mn5@105_d N_OUT4_Mn5@105_g N_VSS_Mn5@105_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@104 N_OUT5_Mn5@104_d N_OUT4_Mn5@104_g N_VSS_Mn5@104_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@105 N_OUT5_Mp5@105_d N_OUT4_Mp5@105_g N_VDD_Mp5@105_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@104 N_OUT5_Mp5@104_d N_OUT4_Mp5@104_g N_VDD_Mp5@104_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@103 N_OUT5_Mn5@103_d N_OUT4_Mn5@103_g N_VSS_Mn5@103_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@102 N_OUT5_Mn5@102_d N_OUT4_Mn5@102_g N_VSS_Mn5@102_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@103 N_OUT5_Mp5@103_d N_OUT4_Mp5@103_g N_VDD_Mp5@103_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@102 N_OUT5_Mp5@102_d N_OUT4_Mp5@102_g N_VDD_Mp5@102_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@101 N_OUT5_Mn5@101_d N_OUT4_Mn5@101_g N_VSS_Mn5@101_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@100 N_OUT5_Mn5@100_d N_OUT4_Mn5@100_g N_VSS_Mn5@100_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@101 N_OUT5_Mp5@101_d N_OUT4_Mp5@101_g N_VDD_Mp5@101_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@100 N_OUT5_Mp5@100_d N_OUT4_Mp5@100_g N_VDD_Mp5@100_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@99 N_OUT5_Mn5@99_d N_OUT4_Mn5@99_g N_VSS_Mn5@99_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@98 N_OUT5_Mn5@98_d N_OUT4_Mn5@98_g N_VSS_Mn5@98_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@99 N_OUT5_Mp5@99_d N_OUT4_Mp5@99_g N_VDD_Mp5@99_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@98 N_OUT5_Mp5@98_d N_OUT4_Mp5@98_g N_VDD_Mp5@98_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3769 N_OUT8_Mn8@3769_d N_OUT7_Mn8@3769_g N_VSS_Mn8@3769_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3768 N_OUT8_Mn8@3768_d N_OUT7_Mn8@3768_g N_VSS_Mn8@3768_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3769 N_OUT8_Mp8@3769_d N_OUT7_Mp8@3769_g N_VDD_Mp8@3769_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3768 N_OUT8_Mp8@3768_d N_OUT7_Mp8@3768_g N_VDD_Mp8@3768_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3767 N_OUT8_Mn8@3767_d N_OUT7_Mn8@3767_g N_VSS_Mn8@3767_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3766 N_OUT8_Mn8@3766_d N_OUT7_Mn8@3766_g N_VSS_Mn8@3766_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3767 N_OUT8_Mp8@3767_d N_OUT7_Mp8@3767_g N_VDD_Mp8@3767_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3766 N_OUT8_Mp8@3766_d N_OUT7_Mp8@3766_g N_VDD_Mp8@3766_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3765 N_OUT8_Mn8@3765_d N_OUT7_Mn8@3765_g N_VSS_Mn8@3765_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3764 N_OUT8_Mn8@3764_d N_OUT7_Mn8@3764_g N_VSS_Mn8@3764_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3765 N_OUT8_Mp8@3765_d N_OUT7_Mp8@3765_g N_VDD_Mp8@3765_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3764 N_OUT8_Mp8@3764_d N_OUT7_Mp8@3764_g N_VDD_Mp8@3764_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3763 N_OUT8_Mn8@3763_d N_OUT7_Mn8@3763_g N_VSS_Mn8@3763_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3762 N_OUT8_Mn8@3762_d N_OUT7_Mn8@3762_g N_VSS_Mn8@3762_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3763 N_OUT8_Mp8@3763_d N_OUT7_Mp8@3763_g N_VDD_Mp8@3763_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3762 N_OUT8_Mp8@3762_d N_OUT7_Mp8@3762_g N_VDD_Mp8@3762_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3761 N_OUT8_Mn8@3761_d N_OUT7_Mn8@3761_g N_VSS_Mn8@3761_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3760 N_OUT8_Mn8@3760_d N_OUT7_Mn8@3760_g N_VSS_Mn8@3760_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3761 N_OUT8_Mp8@3761_d N_OUT7_Mp8@3761_g N_VDD_Mp8@3761_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3760 N_OUT8_Mp8@3760_d N_OUT7_Mp8@3760_g N_VDD_Mp8@3760_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3759 N_OUT8_Mn8@3759_d N_OUT7_Mn8@3759_g N_VSS_Mn8@3759_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3758 N_OUT8_Mn8@3758_d N_OUT7_Mn8@3758_g N_VSS_Mn8@3758_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3759 N_OUT8_Mp8@3759_d N_OUT7_Mp8@3759_g N_VDD_Mp8@3759_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3758 N_OUT8_Mp8@3758_d N_OUT7_Mp8@3758_g N_VDD_Mp8@3758_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3757 N_OUT8_Mn8@3757_d N_OUT7_Mn8@3757_g N_VSS_Mn8@3757_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3756 N_OUT8_Mn8@3756_d N_OUT7_Mn8@3756_g N_VSS_Mn8@3756_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3757 N_OUT8_Mp8@3757_d N_OUT7_Mp8@3757_g N_VDD_Mp8@3757_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3756 N_OUT8_Mp8@3756_d N_OUT7_Mp8@3756_g N_VDD_Mp8@3756_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3755 N_OUT8_Mn8@3755_d N_OUT7_Mn8@3755_g N_VSS_Mn8@3755_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3754 N_OUT8_Mn8@3754_d N_OUT7_Mn8@3754_g N_VSS_Mn8@3754_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3755 N_OUT8_Mp8@3755_d N_OUT7_Mp8@3755_g N_VDD_Mp8@3755_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3754 N_OUT8_Mp8@3754_d N_OUT7_Mp8@3754_g N_VDD_Mp8@3754_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3753 N_OUT8_Mn8@3753_d N_OUT7_Mn8@3753_g N_VSS_Mn8@3753_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3752 N_OUT8_Mn8@3752_d N_OUT7_Mn8@3752_g N_VSS_Mn8@3752_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3753 N_OUT8_Mp8@3753_d N_OUT7_Mp8@3753_g N_VDD_Mp8@3753_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3752 N_OUT8_Mp8@3752_d N_OUT7_Mp8@3752_g N_VDD_Mp8@3752_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3751 N_OUT8_Mn8@3751_d N_OUT7_Mn8@3751_g N_VSS_Mn8@3751_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3750 N_OUT8_Mn8@3750_d N_OUT7_Mn8@3750_g N_VSS_Mn8@3750_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3751 N_OUT8_Mp8@3751_d N_OUT7_Mp8@3751_g N_VDD_Mp8@3751_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3750 N_OUT8_Mp8@3750_d N_OUT7_Mp8@3750_g N_VDD_Mp8@3750_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3749 N_OUT8_Mn8@3749_d N_OUT7_Mn8@3749_g N_VSS_Mn8@3749_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3748 N_OUT8_Mn8@3748_d N_OUT7_Mn8@3748_g N_VSS_Mn8@3748_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3749 N_OUT8_Mp8@3749_d N_OUT7_Mp8@3749_g N_VDD_Mp8@3749_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3748 N_OUT8_Mp8@3748_d N_OUT7_Mp8@3748_g N_VDD_Mp8@3748_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3747 N_OUT8_Mn8@3747_d N_OUT7_Mn8@3747_g N_VSS_Mn8@3747_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3746 N_OUT8_Mn8@3746_d N_OUT7_Mn8@3746_g N_VSS_Mn8@3746_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3747 N_OUT8_Mp8@3747_d N_OUT7_Mp8@3747_g N_VDD_Mp8@3747_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3746 N_OUT8_Mp8@3746_d N_OUT7_Mp8@3746_g N_VDD_Mp8@3746_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@97 N_OUT5_Mn5@97_d N_OUT4_Mn5@97_g N_VSS_Mn5@97_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@96 N_OUT5_Mn5@96_d N_OUT4_Mn5@96_g N_VSS_Mn5@96_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@97 N_OUT5_Mp5@97_d N_OUT4_Mp5@97_g N_VDD_Mp5@97_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@96 N_OUT5_Mp5@96_d N_OUT4_Mp5@96_g N_VDD_Mp5@96_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@95 N_OUT5_Mn5@95_d N_OUT4_Mn5@95_g N_VSS_Mn5@95_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@94 N_OUT5_Mn5@94_d N_OUT4_Mn5@94_g N_VSS_Mn5@94_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@95 N_OUT5_Mp5@95_d N_OUT4_Mp5@95_g N_VDD_Mp5@95_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@94 N_OUT5_Mp5@94_d N_OUT4_Mp5@94_g N_VDD_Mp5@94_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@93 N_OUT5_Mn5@93_d N_OUT4_Mn5@93_g N_VSS_Mn5@93_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@92 N_OUT5_Mn5@92_d N_OUT4_Mn5@92_g N_VSS_Mn5@92_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@93 N_OUT5_Mp5@93_d N_OUT4_Mp5@93_g N_VDD_Mp5@93_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@92 N_OUT5_Mp5@92_d N_OUT4_Mp5@92_g N_VDD_Mp5@92_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@91 N_OUT5_Mn5@91_d N_OUT4_Mn5@91_g N_VSS_Mn5@91_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@90 N_OUT5_Mn5@90_d N_OUT4_Mn5@90_g N_VSS_Mn5@90_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@91 N_OUT5_Mp5@91_d N_OUT4_Mp5@91_g N_VDD_Mp5@91_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@90 N_OUT5_Mp5@90_d N_OUT4_Mp5@90_g N_VDD_Mp5@90_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@89 N_OUT5_Mn5@89_d N_OUT4_Mn5@89_g N_VSS_Mn5@89_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@88 N_OUT5_Mn5@88_d N_OUT4_Mn5@88_g N_VSS_Mn5@88_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@89 N_OUT5_Mp5@89_d N_OUT4_Mp5@89_g N_VDD_Mp5@89_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@88 N_OUT5_Mp5@88_d N_OUT4_Mp5@88_g N_VDD_Mp5@88_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@87 N_OUT5_Mn5@87_d N_OUT4_Mn5@87_g N_VSS_Mn5@87_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@86 N_OUT5_Mn5@86_d N_OUT4_Mn5@86_g N_VSS_Mn5@86_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@87 N_OUT5_Mp5@87_d N_OUT4_Mp5@87_g N_VDD_Mp5@87_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@86 N_OUT5_Mp5@86_d N_OUT4_Mp5@86_g N_VDD_Mp5@86_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@85 N_OUT5_Mn5@85_d N_OUT4_Mn5@85_g N_VSS_Mn5@85_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@84 N_OUT5_Mn5@84_d N_OUT4_Mn5@84_g N_VSS_Mn5@84_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@85 N_OUT5_Mp5@85_d N_OUT4_Mp5@85_g N_VDD_Mp5@85_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@84 N_OUT5_Mp5@84_d N_OUT4_Mp5@84_g N_VDD_Mp5@84_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@83 N_OUT5_Mn5@83_d N_OUT4_Mn5@83_g N_VSS_Mn5@83_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@82 N_OUT5_Mn5@82_d N_OUT4_Mn5@82_g N_VSS_Mn5@82_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@83 N_OUT5_Mp5@83_d N_OUT4_Mp5@83_g N_VDD_Mp5@83_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@82 N_OUT5_Mp5@82_d N_OUT4_Mp5@82_g N_VDD_Mp5@82_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@81 N_OUT5_Mn5@81_d N_OUT4_Mn5@81_g N_VSS_Mn5@81_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@80 N_OUT5_Mn5@80_d N_OUT4_Mn5@80_g N_VSS_Mn5@80_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@81 N_OUT5_Mp5@81_d N_OUT4_Mp5@81_g N_VDD_Mp5@81_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@80 N_OUT5_Mp5@80_d N_OUT4_Mp5@80_g N_VDD_Mp5@80_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@79 N_OUT5_Mn5@79_d N_OUT4_Mn5@79_g N_VSS_Mn5@79_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@78 N_OUT5_Mn5@78_d N_OUT4_Mn5@78_g N_VSS_Mn5@78_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@79 N_OUT5_Mp5@79_d N_OUT4_Mp5@79_g N_VDD_Mp5@79_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@78 N_OUT5_Mp5@78_d N_OUT4_Mp5@78_g N_VDD_Mp5@78_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@77 N_OUT5_Mn5@77_d N_OUT4_Mn5@77_g N_VSS_Mn5@77_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@76 N_OUT5_Mn5@76_d N_OUT4_Mn5@76_g N_VSS_Mn5@76_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@77 N_OUT5_Mp5@77_d N_OUT4_Mp5@77_g N_VDD_Mp5@77_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@76 N_OUT5_Mp5@76_d N_OUT4_Mp5@76_g N_VDD_Mp5@76_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@75 N_OUT5_Mn5@75_d N_OUT4_Mn5@75_g N_VSS_Mn5@75_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@74 N_OUT5_Mn5@74_d N_OUT4_Mn5@74_g N_VSS_Mn5@74_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@75 N_OUT5_Mp5@75_d N_OUT4_Mp5@75_g N_VDD_Mp5@75_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@74 N_OUT5_Mp5@74_d N_OUT4_Mp5@74_g N_VDD_Mp5@74_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@73 N_OUT5_Mn5@73_d N_OUT4_Mn5@73_g N_VSS_Mn5@73_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@72 N_OUT5_Mn5@72_d N_OUT4_Mn5@72_g N_VSS_Mn5@72_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@73 N_OUT5_Mp5@73_d N_OUT4_Mp5@73_g N_VDD_Mp5@73_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@72 N_OUT5_Mp5@72_d N_OUT4_Mp5@72_g N_VDD_Mp5@72_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@71 N_OUT5_Mn5@71_d N_OUT4_Mn5@71_g N_VSS_Mn5@71_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@70 N_OUT5_Mn5@70_d N_OUT4_Mn5@70_g N_VSS_Mn5@70_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@71 N_OUT5_Mp5@71_d N_OUT4_Mp5@71_g N_VDD_Mp5@71_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@70 N_OUT5_Mp5@70_d N_OUT4_Mp5@70_g N_VDD_Mp5@70_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@69 N_OUT5_Mn5@69_d N_OUT4_Mn5@69_g N_VSS_Mn5@69_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@68 N_OUT5_Mn5@68_d N_OUT4_Mn5@68_g N_VSS_Mn5@68_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@69 N_OUT5_Mp5@69_d N_OUT4_Mp5@69_g N_VDD_Mp5@69_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@68 N_OUT5_Mp5@68_d N_OUT4_Mp5@68_g N_VDD_Mp5@68_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@67 N_OUT5_Mn5@67_d N_OUT4_Mn5@67_g N_VSS_Mn5@67_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@66 N_OUT5_Mn5@66_d N_OUT4_Mn5@66_g N_VSS_Mn5@66_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@67 N_OUT5_Mp5@67_d N_OUT4_Mp5@67_g N_VDD_Mp5@67_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@66 N_OUT5_Mp5@66_d N_OUT4_Mp5@66_g N_VDD_Mp5@66_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3745 N_OUT8_Mn8@3745_d N_OUT7_Mn8@3745_g N_VSS_Mn8@3745_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3744 N_OUT8_Mn8@3744_d N_OUT7_Mn8@3744_g N_VSS_Mn8@3744_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3745 N_OUT8_Mp8@3745_d N_OUT7_Mp8@3745_g N_VDD_Mp8@3745_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3744 N_OUT8_Mp8@3744_d N_OUT7_Mp8@3744_g N_VDD_Mp8@3744_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3743 N_OUT8_Mn8@3743_d N_OUT7_Mn8@3743_g N_VSS_Mn8@3743_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3742 N_OUT8_Mn8@3742_d N_OUT7_Mn8@3742_g N_VSS_Mn8@3742_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3743 N_OUT8_Mp8@3743_d N_OUT7_Mp8@3743_g N_VDD_Mp8@3743_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3742 N_OUT8_Mp8@3742_d N_OUT7_Mp8@3742_g N_VDD_Mp8@3742_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3741 N_OUT8_Mn8@3741_d N_OUT7_Mn8@3741_g N_VSS_Mn8@3741_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3740 N_OUT8_Mn8@3740_d N_OUT7_Mn8@3740_g N_VSS_Mn8@3740_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3741 N_OUT8_Mp8@3741_d N_OUT7_Mp8@3741_g N_VDD_Mp8@3741_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3740 N_OUT8_Mp8@3740_d N_OUT7_Mp8@3740_g N_VDD_Mp8@3740_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3739 N_OUT8_Mn8@3739_d N_OUT7_Mn8@3739_g N_VSS_Mn8@3739_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3738 N_OUT8_Mn8@3738_d N_OUT7_Mn8@3738_g N_VSS_Mn8@3738_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3739 N_OUT8_Mp8@3739_d N_OUT7_Mp8@3739_g N_VDD_Mp8@3739_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3738 N_OUT8_Mp8@3738_d N_OUT7_Mp8@3738_g N_VDD_Mp8@3738_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3737 N_OUT8_Mn8@3737_d N_OUT7_Mn8@3737_g N_VSS_Mn8@3737_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3736 N_OUT8_Mn8@3736_d N_OUT7_Mn8@3736_g N_VSS_Mn8@3736_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3737 N_OUT8_Mp8@3737_d N_OUT7_Mp8@3737_g N_VDD_Mp8@3737_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3736 N_OUT8_Mp8@3736_d N_OUT7_Mp8@3736_g N_VDD_Mp8@3736_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3735 N_OUT8_Mn8@3735_d N_OUT7_Mn8@3735_g N_VSS_Mn8@3735_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3734 N_OUT8_Mn8@3734_d N_OUT7_Mn8@3734_g N_VSS_Mn8@3734_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3735 N_OUT8_Mp8@3735_d N_OUT7_Mp8@3735_g N_VDD_Mp8@3735_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3734 N_OUT8_Mp8@3734_d N_OUT7_Mp8@3734_g N_VDD_Mp8@3734_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3733 N_OUT8_Mn8@3733_d N_OUT7_Mn8@3733_g N_VSS_Mn8@3733_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3732 N_OUT8_Mn8@3732_d N_OUT7_Mn8@3732_g N_VSS_Mn8@3732_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3733 N_OUT8_Mp8@3733_d N_OUT7_Mp8@3733_g N_VDD_Mp8@3733_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3732 N_OUT8_Mp8@3732_d N_OUT7_Mp8@3732_g N_VDD_Mp8@3732_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3731 N_OUT8_Mn8@3731_d N_OUT7_Mn8@3731_g N_VSS_Mn8@3731_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3730 N_OUT8_Mn8@3730_d N_OUT7_Mn8@3730_g N_VSS_Mn8@3730_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3731 N_OUT8_Mp8@3731_d N_OUT7_Mp8@3731_g N_VDD_Mp8@3731_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3730 N_OUT8_Mp8@3730_d N_OUT7_Mp8@3730_g N_VDD_Mp8@3730_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3729 N_OUT8_Mn8@3729_d N_OUT7_Mn8@3729_g N_VSS_Mn8@3729_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3728 N_OUT8_Mn8@3728_d N_OUT7_Mn8@3728_g N_VSS_Mn8@3728_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3729 N_OUT8_Mp8@3729_d N_OUT7_Mp8@3729_g N_VDD_Mp8@3729_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3728 N_OUT8_Mp8@3728_d N_OUT7_Mp8@3728_g N_VDD_Mp8@3728_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3727 N_OUT8_Mn8@3727_d N_OUT7_Mn8@3727_g N_VSS_Mn8@3727_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3726 N_OUT8_Mn8@3726_d N_OUT7_Mn8@3726_g N_VSS_Mn8@3726_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3727 N_OUT8_Mp8@3727_d N_OUT7_Mp8@3727_g N_VDD_Mp8@3727_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3726 N_OUT8_Mp8@3726_d N_OUT7_Mp8@3726_g N_VDD_Mp8@3726_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3725 N_OUT8_Mn8@3725_d N_OUT7_Mn8@3725_g N_VSS_Mn8@3725_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3724 N_OUT8_Mn8@3724_d N_OUT7_Mn8@3724_g N_VSS_Mn8@3724_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3725 N_OUT8_Mp8@3725_d N_OUT7_Mp8@3725_g N_VDD_Mp8@3725_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3724 N_OUT8_Mp8@3724_d N_OUT7_Mp8@3724_g N_VDD_Mp8@3724_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3723 N_OUT8_Mn8@3723_d N_OUT7_Mn8@3723_g N_VSS_Mn8@3723_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3722 N_OUT8_Mn8@3722_d N_OUT7_Mn8@3722_g N_VSS_Mn8@3722_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3723 N_OUT8_Mp8@3723_d N_OUT7_Mp8@3723_g N_VDD_Mp8@3723_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3722 N_OUT8_Mp8@3722_d N_OUT7_Mp8@3722_g N_VDD_Mp8@3722_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3721 N_OUT8_Mn8@3721_d N_OUT7_Mn8@3721_g N_VSS_Mn8@3721_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3720 N_OUT8_Mn8@3720_d N_OUT7_Mn8@3720_g N_VSS_Mn8@3720_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3721 N_OUT8_Mp8@3721_d N_OUT7_Mp8@3721_g N_VDD_Mp8@3721_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3720 N_OUT8_Mp8@3720_d N_OUT7_Mp8@3720_g N_VDD_Mp8@3720_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3719 N_OUT8_Mn8@3719_d N_OUT7_Mn8@3719_g N_VSS_Mn8@3719_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3718 N_OUT8_Mn8@3718_d N_OUT7_Mn8@3718_g N_VSS_Mn8@3718_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3719 N_OUT8_Mp8@3719_d N_OUT7_Mp8@3719_g N_VDD_Mp8@3719_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3718 N_OUT8_Mp8@3718_d N_OUT7_Mp8@3718_g N_VDD_Mp8@3718_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3717 N_OUT8_Mn8@3717_d N_OUT7_Mn8@3717_g N_VSS_Mn8@3717_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3716 N_OUT8_Mn8@3716_d N_OUT7_Mn8@3716_g N_VSS_Mn8@3716_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3717 N_OUT8_Mp8@3717_d N_OUT7_Mp8@3717_g N_VDD_Mp8@3717_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3716 N_OUT8_Mp8@3716_d N_OUT7_Mp8@3716_g N_VDD_Mp8@3716_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3715 N_OUT8_Mn8@3715_d N_OUT7_Mn8@3715_g N_VSS_Mn8@3715_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3714 N_OUT8_Mn8@3714_d N_OUT7_Mn8@3714_g N_VSS_Mn8@3714_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3715 N_OUT8_Mp8@3715_d N_OUT7_Mp8@3715_g N_VDD_Mp8@3715_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3714 N_OUT8_Mp8@3714_d N_OUT7_Mp8@3714_g N_VDD_Mp8@3714_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@65 N_OUT5_Mn5@65_d N_OUT4_Mn5@65_g N_VSS_Mn5@65_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@64 N_OUT5_Mn5@64_d N_OUT4_Mn5@64_g N_VSS_Mn5@64_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@65 N_OUT5_Mp5@65_d N_OUT4_Mp5@65_g N_VDD_Mp5@65_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@64 N_OUT5_Mp5@64_d N_OUT4_Mp5@64_g N_VDD_Mp5@64_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@63 N_OUT5_Mn5@63_d N_OUT4_Mn5@63_g N_VSS_Mn5@63_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@62 N_OUT5_Mn5@62_d N_OUT4_Mn5@62_g N_VSS_Mn5@62_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@63 N_OUT5_Mp5@63_d N_OUT4_Mp5@63_g N_VDD_Mp5@63_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@62 N_OUT5_Mp5@62_d N_OUT4_Mp5@62_g N_VDD_Mp5@62_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@61 N_OUT5_Mn5@61_d N_OUT4_Mn5@61_g N_VSS_Mn5@61_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@60 N_OUT5_Mn5@60_d N_OUT4_Mn5@60_g N_VSS_Mn5@60_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@61 N_OUT5_Mp5@61_d N_OUT4_Mp5@61_g N_VDD_Mp5@61_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@60 N_OUT5_Mp5@60_d N_OUT4_Mp5@60_g N_VDD_Mp5@60_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@59 N_OUT5_Mn5@59_d N_OUT4_Mn5@59_g N_VSS_Mn5@59_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@58 N_OUT5_Mn5@58_d N_OUT4_Mn5@58_g N_VSS_Mn5@58_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@59 N_OUT5_Mp5@59_d N_OUT4_Mp5@59_g N_VDD_Mp5@59_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@58 N_OUT5_Mp5@58_d N_OUT4_Mp5@58_g N_VDD_Mp5@58_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@57 N_OUT5_Mn5@57_d N_OUT4_Mn5@57_g N_VSS_Mn5@57_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@56 N_OUT5_Mn5@56_d N_OUT4_Mn5@56_g N_VSS_Mn5@56_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@57 N_OUT5_Mp5@57_d N_OUT4_Mp5@57_g N_VDD_Mp5@57_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@56 N_OUT5_Mp5@56_d N_OUT4_Mp5@56_g N_VDD_Mp5@56_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@55 N_OUT5_Mn5@55_d N_OUT4_Mn5@55_g N_VSS_Mn5@55_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@54 N_OUT5_Mn5@54_d N_OUT4_Mn5@54_g N_VSS_Mn5@54_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@55 N_OUT5_Mp5@55_d N_OUT4_Mp5@55_g N_VDD_Mp5@55_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@54 N_OUT5_Mp5@54_d N_OUT4_Mp5@54_g N_VDD_Mp5@54_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@53 N_OUT5_Mn5@53_d N_OUT4_Mn5@53_g N_VSS_Mn5@53_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@52 N_OUT5_Mn5@52_d N_OUT4_Mn5@52_g N_VSS_Mn5@52_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@53 N_OUT5_Mp5@53_d N_OUT4_Mp5@53_g N_VDD_Mp5@53_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@52 N_OUT5_Mp5@52_d N_OUT4_Mp5@52_g N_VDD_Mp5@52_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@51 N_OUT5_Mn5@51_d N_OUT4_Mn5@51_g N_VSS_Mn5@51_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@50 N_OUT5_Mn5@50_d N_OUT4_Mn5@50_g N_VSS_Mn5@50_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@51 N_OUT5_Mp5@51_d N_OUT4_Mp5@51_g N_VDD_Mp5@51_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@50 N_OUT5_Mp5@50_d N_OUT4_Mp5@50_g N_VDD_Mp5@50_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@49 N_OUT5_Mn5@49_d N_OUT4_Mn5@49_g N_VSS_Mn5@49_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@48 N_OUT5_Mn5@48_d N_OUT4_Mn5@48_g N_VSS_Mn5@48_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@49 N_OUT5_Mp5@49_d N_OUT4_Mp5@49_g N_VDD_Mp5@49_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@48 N_OUT5_Mp5@48_d N_OUT4_Mp5@48_g N_VDD_Mp5@48_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@47 N_OUT5_Mn5@47_d N_OUT4_Mn5@47_g N_VSS_Mn5@47_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@46 N_OUT5_Mn5@46_d N_OUT4_Mn5@46_g N_VSS_Mn5@46_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@47 N_OUT5_Mp5@47_d N_OUT4_Mp5@47_g N_VDD_Mp5@47_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@46 N_OUT5_Mp5@46_d N_OUT4_Mp5@46_g N_VDD_Mp5@46_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@45 N_OUT5_Mn5@45_d N_OUT4_Mn5@45_g N_VSS_Mn5@45_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@44 N_OUT5_Mn5@44_d N_OUT4_Mn5@44_g N_VSS_Mn5@44_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@45 N_OUT5_Mp5@45_d N_OUT4_Mp5@45_g N_VDD_Mp5@45_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@44 N_OUT5_Mp5@44_d N_OUT4_Mp5@44_g N_VDD_Mp5@44_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@43 N_OUT5_Mn5@43_d N_OUT4_Mn5@43_g N_VSS_Mn5@43_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@42 N_OUT5_Mn5@42_d N_OUT4_Mn5@42_g N_VSS_Mn5@42_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@43 N_OUT5_Mp5@43_d N_OUT4_Mp5@43_g N_VDD_Mp5@43_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@42 N_OUT5_Mp5@42_d N_OUT4_Mp5@42_g N_VDD_Mp5@42_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@41 N_OUT5_Mn5@41_d N_OUT4_Mn5@41_g N_VSS_Mn5@41_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@40 N_OUT5_Mn5@40_d N_OUT4_Mn5@40_g N_VSS_Mn5@40_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@41 N_OUT5_Mp5@41_d N_OUT4_Mp5@41_g N_VDD_Mp5@41_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@40 N_OUT5_Mp5@40_d N_OUT4_Mp5@40_g N_VDD_Mp5@40_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@39 N_OUT5_Mn5@39_d N_OUT4_Mn5@39_g N_VSS_Mn5@39_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@38 N_OUT5_Mn5@38_d N_OUT4_Mn5@38_g N_VSS_Mn5@38_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@39 N_OUT5_Mp5@39_d N_OUT4_Mp5@39_g N_VDD_Mp5@39_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@38 N_OUT5_Mp5@38_d N_OUT4_Mp5@38_g N_VDD_Mp5@38_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@37 N_OUT5_Mn5@37_d N_OUT4_Mn5@37_g N_VSS_Mn5@37_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@36 N_OUT5_Mn5@36_d N_OUT4_Mn5@36_g N_VSS_Mn5@36_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@37 N_OUT5_Mp5@37_d N_OUT4_Mp5@37_g N_VDD_Mp5@37_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@36 N_OUT5_Mp5@36_d N_OUT4_Mp5@36_g N_VDD_Mp5@36_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@35 N_OUT5_Mn5@35_d N_OUT4_Mn5@35_g N_VSS_Mn5@35_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@34 N_OUT5_Mn5@34_d N_OUT4_Mn5@34_g N_VSS_Mn5@34_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@35 N_OUT5_Mp5@35_d N_OUT4_Mp5@35_g N_VDD_Mp5@35_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@34 N_OUT5_Mp5@34_d N_OUT4_Mp5@34_g N_VDD_Mp5@34_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@33 N_OUT5_Mn5@33_d N_OUT4_Mn5@33_g N_VSS_Mn5@33_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@32 N_OUT5_Mn5@32_d N_OUT4_Mn5@32_g N_VSS_Mn5@32_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@33 N_OUT5_Mp5@33_d N_OUT4_Mp5@33_g N_VDD_Mp5@33_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@32 N_OUT5_Mp5@32_d N_OUT4_Mp5@32_g N_VDD_Mp5@32_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@31 N_OUT5_Mn5@31_d N_OUT4_Mn5@31_g N_VSS_Mn5@31_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@30 N_OUT5_Mn5@30_d N_OUT4_Mn5@30_g N_VSS_Mn5@30_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@31 N_OUT5_Mp5@31_d N_OUT4_Mp5@31_g N_VDD_Mp5@31_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@30 N_OUT5_Mp5@30_d N_OUT4_Mp5@30_g N_VDD_Mp5@30_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@29 N_OUT5_Mn5@29_d N_OUT4_Mn5@29_g N_VSS_Mn5@29_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@28 N_OUT5_Mn5@28_d N_OUT4_Mn5@28_g N_VSS_Mn5@28_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@29 N_OUT5_Mp5@29_d N_OUT4_Mp5@29_g N_VDD_Mp5@29_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@28 N_OUT5_Mp5@28_d N_OUT4_Mp5@28_g N_VDD_Mp5@28_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@27 N_OUT5_Mn5@27_d N_OUT4_Mn5@27_g N_VSS_Mn5@27_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@26 N_OUT5_Mn5@26_d N_OUT4_Mn5@26_g N_VSS_Mn5@26_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@27 N_OUT5_Mp5@27_d N_OUT4_Mp5@27_g N_VDD_Mp5@27_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@26 N_OUT5_Mp5@26_d N_OUT4_Mp5@26_g N_VDD_Mp5@26_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@25 N_OUT5_Mn5@25_d N_OUT4_Mn5@25_g N_VSS_Mn5@25_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@24 N_OUT5_Mn5@24_d N_OUT4_Mn5@24_g N_VSS_Mn5@24_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@25 N_OUT5_Mp5@25_d N_OUT4_Mp5@25_g N_VDD_Mp5@25_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@24 N_OUT5_Mp5@24_d N_OUT4_Mp5@24_g N_VDD_Mp5@24_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@23 N_OUT5_Mn5@23_d N_OUT4_Mn5@23_g N_VSS_Mn5@23_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@22 N_OUT5_Mn5@22_d N_OUT4_Mn5@22_g N_VSS_Mn5@22_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@23 N_OUT5_Mp5@23_d N_OUT4_Mp5@23_g N_VDD_Mp5@23_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@22 N_OUT5_Mp5@22_d N_OUT4_Mp5@22_g N_VDD_Mp5@22_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@21 N_OUT5_Mn5@21_d N_OUT4_Mn5@21_g N_VSS_Mn5@21_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@20 N_OUT5_Mn5@20_d N_OUT4_Mn5@20_g N_VSS_Mn5@20_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@21 N_OUT5_Mp5@21_d N_OUT4_Mp5@21_g N_VDD_Mp5@21_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@20 N_OUT5_Mp5@20_d N_OUT4_Mp5@20_g N_VDD_Mp5@20_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@19 N_OUT5_Mn5@19_d N_OUT4_Mn5@19_g N_VSS_Mn5@19_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@18 N_OUT5_Mn5@18_d N_OUT4_Mn5@18_g N_VSS_Mn5@18_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@19 N_OUT5_Mp5@19_d N_OUT4_Mp5@19_g N_VDD_Mp5@19_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@18 N_OUT5_Mp5@18_d N_OUT4_Mp5@18_g N_VDD_Mp5@18_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@17 N_OUT5_Mn5@17_d N_OUT4_Mn5@17_g N_VSS_Mn5@17_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@16 N_OUT5_Mn5@16_d N_OUT4_Mn5@16_g N_VSS_Mn5@16_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@17 N_OUT5_Mp5@17_d N_OUT4_Mp5@17_g N_VDD_Mp5@17_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@16 N_OUT5_Mp5@16_d N_OUT4_Mp5@16_g N_VDD_Mp5@16_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@15 N_OUT5_Mn5@15_d N_OUT4_Mn5@15_g N_VSS_Mn5@15_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@14 N_OUT5_Mn5@14_d N_OUT4_Mn5@14_g N_VSS_Mn5@14_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@15 N_OUT5_Mp5@15_d N_OUT4_Mp5@15_g N_VDD_Mp5@15_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@14 N_OUT5_Mp5@14_d N_OUT4_Mp5@14_g N_VDD_Mp5@14_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@13 N_OUT5_Mn5@13_d N_OUT4_Mn5@13_g N_VSS_Mn5@13_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@12 N_OUT5_Mn5@12_d N_OUT4_Mn5@12_g N_VSS_Mn5@12_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@13 N_OUT5_Mp5@13_d N_OUT4_Mp5@13_g N_VDD_Mp5@13_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@12 N_OUT5_Mp5@12_d N_OUT4_Mp5@12_g N_VDD_Mp5@12_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@11 N_OUT5_Mn5@11_d N_OUT4_Mn5@11_g N_VSS_Mn5@11_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@10 N_OUT5_Mn5@10_d N_OUT4_Mn5@10_g N_VSS_Mn5@10_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@11 N_OUT5_Mp5@11_d N_OUT4_Mp5@11_g N_VDD_Mp5@11_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@10 N_OUT5_Mp5@10_d N_OUT4_Mp5@10_g N_VDD_Mp5@10_s N_VDD_Mp5@105_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@9 N_OUT5_Mn5@9_d N_OUT4_Mn5@9_g N_VSS_Mn5@9_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@8 N_OUT5_Mn5@8_d N_OUT4_Mn5@8_g N_VSS_Mn5@8_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@9 N_OUT5_Mp5@9_d N_OUT4_Mp5@9_g N_VDD_Mp5@9_s N_VDD_Mp5@105_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@8 N_OUT5_Mp5@8_d N_OUT4_Mp5@8_g N_VDD_Mp5@8_s N_VDD_Mp5@105_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@7 N_OUT5_Mn5@7_d N_OUT4_Mn5@7_g N_VSS_Mn5@7_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@6 N_OUT5_Mn5@6_d N_OUT4_Mn5@6_g N_VSS_Mn5@6_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@7 N_OUT5_Mp5@7_d N_OUT4_Mp5@7_g N_VDD_Mp5@7_s N_VDD_Mp5@105_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@6 N_OUT5_Mp5@6_d N_OUT4_Mp5@6_g N_VDD_Mp5@6_s N_VDD_Mp5@105_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@5 N_OUT5_Mn5@5_d N_OUT4_Mn5@5_g N_VSS_Mn5@5_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@4 N_OUT5_Mn5@4_d N_OUT4_Mn5@4_g N_VSS_Mn5@4_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@5 N_OUT5_Mp5@5_d N_OUT4_Mp5@5_g N_VDD_Mp5@5_s N_VDD_Mp5@105_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@4 N_OUT5_Mp5@4_d N_OUT4_Mp5@4_g N_VDD_Mp5@4_s N_VDD_Mp5@105_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn5@3 N_OUT5_Mn5@3_d N_OUT4_Mn5@3_g N_VSS_Mn5@3_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn5@2 N_OUT5_Mn5@2_d N_OUT4_Mn5@2_g N_VSS_Mn5@2_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp5@3 N_OUT5_Mp5@3_d N_OUT4_Mp5@3_g N_VDD_Mp5@3_s N_VDD_Mp5@105_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp5@2 N_OUT5_Mp5@2_d N_OUT4_Mp5@2_g N_VDD_Mp5@2_s N_VDD_Mp5@105_b P_18 L=1.8e-07
+ W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1153 N_OUT7_Mn7@1153_d N_OUT6_Mn7@1153_g N_VSS_Mn7@1153_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1152 N_OUT7_Mn7@1152_d N_OUT6_Mn7@1152_g N_VSS_Mn7@1152_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1153 N_OUT7_Mp7@1153_d N_OUT6_Mp7@1153_g N_VDD_Mp7@1153_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1152 N_OUT7_Mp7@1152_d N_OUT6_Mp7@1152_g N_VDD_Mp7@1152_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1151 N_OUT7_Mn7@1151_d N_OUT6_Mn7@1151_g N_VSS_Mn7@1151_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1150 N_OUT7_Mn7@1150_d N_OUT6_Mn7@1150_g N_VSS_Mn7@1150_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1151 N_OUT7_Mp7@1151_d N_OUT6_Mp7@1151_g N_VDD_Mp7@1151_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1150 N_OUT7_Mp7@1150_d N_OUT6_Mp7@1150_g N_VDD_Mp7@1150_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1149 N_OUT7_Mn7@1149_d N_OUT6_Mn7@1149_g N_VSS_Mn7@1149_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1148 N_OUT7_Mn7@1148_d N_OUT6_Mn7@1148_g N_VSS_Mn7@1148_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1149 N_OUT7_Mp7@1149_d N_OUT6_Mp7@1149_g N_VDD_Mp7@1149_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1148 N_OUT7_Mp7@1148_d N_OUT6_Mp7@1148_g N_VDD_Mp7@1148_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1147 N_OUT7_Mn7@1147_d N_OUT6_Mn7@1147_g N_VSS_Mn7@1147_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1146 N_OUT7_Mn7@1146_d N_OUT6_Mn7@1146_g N_VSS_Mn7@1146_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1147 N_OUT7_Mp7@1147_d N_OUT6_Mp7@1147_g N_VDD_Mp7@1147_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1146 N_OUT7_Mp7@1146_d N_OUT6_Mp7@1146_g N_VDD_Mp7@1146_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1145 N_OUT7_Mn7@1145_d N_OUT6_Mn7@1145_g N_VSS_Mn7@1145_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1144 N_OUT7_Mn7@1144_d N_OUT6_Mn7@1144_g N_VSS_Mn7@1144_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1145 N_OUT7_Mp7@1145_d N_OUT6_Mp7@1145_g N_VDD_Mp7@1145_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1144 N_OUT7_Mp7@1144_d N_OUT6_Mp7@1144_g N_VDD_Mp7@1144_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1143 N_OUT7_Mn7@1143_d N_OUT6_Mn7@1143_g N_VSS_Mn7@1143_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1142 N_OUT7_Mn7@1142_d N_OUT6_Mn7@1142_g N_VSS_Mn7@1142_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1143 N_OUT7_Mp7@1143_d N_OUT6_Mp7@1143_g N_VDD_Mp7@1143_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1142 N_OUT7_Mp7@1142_d N_OUT6_Mp7@1142_g N_VDD_Mp7@1142_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1141 N_OUT7_Mn7@1141_d N_OUT6_Mn7@1141_g N_VSS_Mn7@1141_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1140 N_OUT7_Mn7@1140_d N_OUT6_Mn7@1140_g N_VSS_Mn7@1140_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1141 N_OUT7_Mp7@1141_d N_OUT6_Mp7@1141_g N_VDD_Mp7@1141_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1140 N_OUT7_Mp7@1140_d N_OUT6_Mp7@1140_g N_VDD_Mp7@1140_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1139 N_OUT7_Mn7@1139_d N_OUT6_Mn7@1139_g N_VSS_Mn7@1139_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1138 N_OUT7_Mn7@1138_d N_OUT6_Mn7@1138_g N_VSS_Mn7@1138_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1139 N_OUT7_Mp7@1139_d N_OUT6_Mp7@1139_g N_VDD_Mp7@1139_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1138 N_OUT7_Mp7@1138_d N_OUT6_Mp7@1138_g N_VDD_Mp7@1138_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1137 N_OUT7_Mn7@1137_d N_OUT6_Mn7@1137_g N_VSS_Mn7@1137_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1136 N_OUT7_Mn7@1136_d N_OUT6_Mn7@1136_g N_VSS_Mn7@1136_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1137 N_OUT7_Mp7@1137_d N_OUT6_Mp7@1137_g N_VDD_Mp7@1137_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1136 N_OUT7_Mp7@1136_d N_OUT6_Mp7@1136_g N_VDD_Mp7@1136_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1135 N_OUT7_Mn7@1135_d N_OUT6_Mn7@1135_g N_VSS_Mn7@1135_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1134 N_OUT7_Mn7@1134_d N_OUT6_Mn7@1134_g N_VSS_Mn7@1134_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1135 N_OUT7_Mp7@1135_d N_OUT6_Mp7@1135_g N_VDD_Mp7@1135_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1134 N_OUT7_Mp7@1134_d N_OUT6_Mp7@1134_g N_VDD_Mp7@1134_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1133 N_OUT7_Mn7@1133_d N_OUT6_Mn7@1133_g N_VSS_Mn7@1133_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1132 N_OUT7_Mn7@1132_d N_OUT6_Mn7@1132_g N_VSS_Mn7@1132_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1133 N_OUT7_Mp7@1133_d N_OUT6_Mp7@1133_g N_VDD_Mp7@1133_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1132 N_OUT7_Mp7@1132_d N_OUT6_Mp7@1132_g N_VDD_Mp7@1132_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1131 N_OUT7_Mn7@1131_d N_OUT6_Mn7@1131_g N_VSS_Mn7@1131_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1130 N_OUT7_Mn7@1130_d N_OUT6_Mn7@1130_g N_VSS_Mn7@1130_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1131 N_OUT7_Mp7@1131_d N_OUT6_Mp7@1131_g N_VDD_Mp7@1131_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1130 N_OUT7_Mp7@1130_d N_OUT6_Mp7@1130_g N_VDD_Mp7@1130_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1129 N_OUT7_Mn7@1129_d N_OUT6_Mn7@1129_g N_VSS_Mn7@1129_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1128 N_OUT7_Mn7@1128_d N_OUT6_Mn7@1128_g N_VSS_Mn7@1128_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1129 N_OUT7_Mp7@1129_d N_OUT6_Mp7@1129_g N_VDD_Mp7@1129_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1128 N_OUT7_Mp7@1128_d N_OUT6_Mp7@1128_g N_VDD_Mp7@1128_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1127 N_OUT7_Mn7@1127_d N_OUT6_Mn7@1127_g N_VSS_Mn7@1127_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1126 N_OUT7_Mn7@1126_d N_OUT6_Mn7@1126_g N_VSS_Mn7@1126_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1127 N_OUT7_Mp7@1127_d N_OUT6_Mp7@1127_g N_VDD_Mp7@1127_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1126 N_OUT7_Mp7@1126_d N_OUT6_Mp7@1126_g N_VDD_Mp7@1126_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1125 N_OUT7_Mn7@1125_d N_OUT6_Mn7@1125_g N_VSS_Mn7@1125_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1124 N_OUT7_Mn7@1124_d N_OUT6_Mn7@1124_g N_VSS_Mn7@1124_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1125 N_OUT7_Mp7@1125_d N_OUT6_Mp7@1125_g N_VDD_Mp7@1125_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1124 N_OUT7_Mp7@1124_d N_OUT6_Mp7@1124_g N_VDD_Mp7@1124_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1123 N_OUT7_Mn7@1123_d N_OUT6_Mn7@1123_g N_VSS_Mn7@1123_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1122 N_OUT7_Mn7@1122_d N_OUT6_Mn7@1122_g N_VSS_Mn7@1122_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1123 N_OUT7_Mp7@1123_d N_OUT6_Mp7@1123_g N_VDD_Mp7@1123_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1122 N_OUT7_Mp7@1122_d N_OUT6_Mp7@1122_g N_VDD_Mp7@1122_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1121 N_OUT7_Mn7@1121_d N_OUT6_Mn7@1121_g N_VSS_Mn7@1121_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1120 N_OUT7_Mn7@1120_d N_OUT6_Mn7@1120_g N_VSS_Mn7@1120_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1121 N_OUT7_Mp7@1121_d N_OUT6_Mp7@1121_g N_VDD_Mp7@1121_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1120 N_OUT7_Mp7@1120_d N_OUT6_Mp7@1120_g N_VDD_Mp7@1120_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1119 N_OUT7_Mn7@1119_d N_OUT6_Mn7@1119_g N_VSS_Mn7@1119_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1118 N_OUT7_Mn7@1118_d N_OUT6_Mn7@1118_g N_VSS_Mn7@1118_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1119 N_OUT7_Mp7@1119_d N_OUT6_Mp7@1119_g N_VDD_Mp7@1119_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1118 N_OUT7_Mp7@1118_d N_OUT6_Mp7@1118_g N_VDD_Mp7@1118_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1117 N_OUT7_Mn7@1117_d N_OUT6_Mn7@1117_g N_VSS_Mn7@1117_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1116 N_OUT7_Mn7@1116_d N_OUT6_Mn7@1116_g N_VSS_Mn7@1116_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1117 N_OUT7_Mp7@1117_d N_OUT6_Mp7@1117_g N_VDD_Mp7@1117_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1116 N_OUT7_Mp7@1116_d N_OUT6_Mp7@1116_g N_VDD_Mp7@1116_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1115 N_OUT7_Mn7@1115_d N_OUT6_Mn7@1115_g N_VSS_Mn7@1115_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1114 N_OUT7_Mn7@1114_d N_OUT6_Mn7@1114_g N_VSS_Mn7@1114_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1115 N_OUT7_Mp7@1115_d N_OUT6_Mp7@1115_g N_VDD_Mp7@1115_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1114 N_OUT7_Mp7@1114_d N_OUT6_Mp7@1114_g N_VDD_Mp7@1114_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1113 N_OUT7_Mn7@1113_d N_OUT6_Mn7@1113_g N_VSS_Mn7@1113_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1112 N_OUT7_Mn7@1112_d N_OUT6_Mn7@1112_g N_VSS_Mn7@1112_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1113 N_OUT7_Mp7@1113_d N_OUT6_Mp7@1113_g N_VDD_Mp7@1113_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1112 N_OUT7_Mp7@1112_d N_OUT6_Mp7@1112_g N_VDD_Mp7@1112_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1111 N_OUT7_Mn7@1111_d N_OUT6_Mn7@1111_g N_VSS_Mn7@1111_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1110 N_OUT7_Mn7@1110_d N_OUT6_Mn7@1110_g N_VSS_Mn7@1110_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1111 N_OUT7_Mp7@1111_d N_OUT6_Mp7@1111_g N_VDD_Mp7@1111_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1110 N_OUT7_Mp7@1110_d N_OUT6_Mp7@1110_g N_VDD_Mp7@1110_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1109 N_OUT7_Mn7@1109_d N_OUT6_Mn7@1109_g N_VSS_Mn7@1109_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1108 N_OUT7_Mn7@1108_d N_OUT6_Mn7@1108_g N_VSS_Mn7@1108_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1109 N_OUT7_Mp7@1109_d N_OUT6_Mp7@1109_g N_VDD_Mp7@1109_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1108 N_OUT7_Mp7@1108_d N_OUT6_Mp7@1108_g N_VDD_Mp7@1108_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1107 N_OUT7_Mn7@1107_d N_OUT6_Mn7@1107_g N_VSS_Mn7@1107_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1106 N_OUT7_Mn7@1106_d N_OUT6_Mn7@1106_g N_VSS_Mn7@1106_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1107 N_OUT7_Mp7@1107_d N_OUT6_Mp7@1107_g N_VDD_Mp7@1107_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1106 N_OUT7_Mp7@1106_d N_OUT6_Mp7@1106_g N_VDD_Mp7@1106_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1105 N_OUT7_Mn7@1105_d N_OUT6_Mn7@1105_g N_VSS_Mn7@1105_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1104 N_OUT7_Mn7@1104_d N_OUT6_Mn7@1104_g N_VSS_Mn7@1104_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1105 N_OUT7_Mp7@1105_d N_OUT6_Mp7@1105_g N_VDD_Mp7@1105_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1104 N_OUT7_Mp7@1104_d N_OUT6_Mp7@1104_g N_VDD_Mp7@1104_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1103 N_OUT7_Mn7@1103_d N_OUT6_Mn7@1103_g N_VSS_Mn7@1103_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1102 N_OUT7_Mn7@1102_d N_OUT6_Mn7@1102_g N_VSS_Mn7@1102_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1103 N_OUT7_Mp7@1103_d N_OUT6_Mp7@1103_g N_VDD_Mp7@1103_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1102 N_OUT7_Mp7@1102_d N_OUT6_Mp7@1102_g N_VDD_Mp7@1102_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1101 N_OUT7_Mn7@1101_d N_OUT6_Mn7@1101_g N_VSS_Mn7@1101_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1100 N_OUT7_Mn7@1100_d N_OUT6_Mn7@1100_g N_VSS_Mn7@1100_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1101 N_OUT7_Mp7@1101_d N_OUT6_Mp7@1101_g N_VDD_Mp7@1101_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1100 N_OUT7_Mp7@1100_d N_OUT6_Mp7@1100_g N_VDD_Mp7@1100_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1099 N_OUT7_Mn7@1099_d N_OUT6_Mn7@1099_g N_VSS_Mn7@1099_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1098 N_OUT7_Mn7@1098_d N_OUT6_Mn7@1098_g N_VSS_Mn7@1098_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1099 N_OUT7_Mp7@1099_d N_OUT6_Mp7@1099_g N_VDD_Mp7@1099_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1098 N_OUT7_Mp7@1098_d N_OUT6_Mp7@1098_g N_VDD_Mp7@1098_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1097 N_OUT7_Mn7@1097_d N_OUT6_Mn7@1097_g N_VSS_Mn7@1097_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1096 N_OUT7_Mn7@1096_d N_OUT6_Mn7@1096_g N_VSS_Mn7@1096_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1097 N_OUT7_Mp7@1097_d N_OUT6_Mp7@1097_g N_VDD_Mp7@1097_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1096 N_OUT7_Mp7@1096_d N_OUT6_Mp7@1096_g N_VDD_Mp7@1096_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1095 N_OUT7_Mn7@1095_d N_OUT6_Mn7@1095_g N_VSS_Mn7@1095_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1094 N_OUT7_Mn7@1094_d N_OUT6_Mn7@1094_g N_VSS_Mn7@1094_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1095 N_OUT7_Mp7@1095_d N_OUT6_Mp7@1095_g N_VDD_Mp7@1095_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1094 N_OUT7_Mp7@1094_d N_OUT6_Mp7@1094_g N_VDD_Mp7@1094_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1093 N_OUT7_Mn7@1093_d N_OUT6_Mn7@1093_g N_VSS_Mn7@1093_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1092 N_OUT7_Mn7@1092_d N_OUT6_Mn7@1092_g N_VSS_Mn7@1092_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1093 N_OUT7_Mp7@1093_d N_OUT6_Mp7@1093_g N_VDD_Mp7@1093_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1092 N_OUT7_Mp7@1092_d N_OUT6_Mp7@1092_g N_VDD_Mp7@1092_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1091 N_OUT7_Mn7@1091_d N_OUT6_Mn7@1091_g N_VSS_Mn7@1091_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1090 N_OUT7_Mn7@1090_d N_OUT6_Mn7@1090_g N_VSS_Mn7@1090_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1091 N_OUT7_Mp7@1091_d N_OUT6_Mp7@1091_g N_VDD_Mp7@1091_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1090 N_OUT7_Mp7@1090_d N_OUT6_Mp7@1090_g N_VDD_Mp7@1090_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1089 N_OUT7_Mn7@1089_d N_OUT6_Mn7@1089_g N_VSS_Mn7@1089_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1088 N_OUT7_Mn7@1088_d N_OUT6_Mn7@1088_g N_VSS_Mn7@1088_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1089 N_OUT7_Mp7@1089_d N_OUT6_Mp7@1089_g N_VDD_Mp7@1089_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1088 N_OUT7_Mp7@1088_d N_OUT6_Mp7@1088_g N_VDD_Mp7@1088_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1087 N_OUT7_Mn7@1087_d N_OUT6_Mn7@1087_g N_VSS_Mn7@1087_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1086 N_OUT7_Mn7@1086_d N_OUT6_Mn7@1086_g N_VSS_Mn7@1086_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1087 N_OUT7_Mp7@1087_d N_OUT6_Mp7@1087_g N_VDD_Mp7@1087_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1086 N_OUT7_Mp7@1086_d N_OUT6_Mp7@1086_g N_VDD_Mp7@1086_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1085 N_OUT7_Mn7@1085_d N_OUT6_Mn7@1085_g N_VSS_Mn7@1085_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1084 N_OUT7_Mn7@1084_d N_OUT6_Mn7@1084_g N_VSS_Mn7@1084_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1085 N_OUT7_Mp7@1085_d N_OUT6_Mp7@1085_g N_VDD_Mp7@1085_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1084 N_OUT7_Mp7@1084_d N_OUT6_Mp7@1084_g N_VDD_Mp7@1084_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1083 N_OUT7_Mn7@1083_d N_OUT6_Mn7@1083_g N_VSS_Mn7@1083_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1082 N_OUT7_Mn7@1082_d N_OUT6_Mn7@1082_g N_VSS_Mn7@1082_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1083 N_OUT7_Mp7@1083_d N_OUT6_Mp7@1083_g N_VDD_Mp7@1083_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1082 N_OUT7_Mp7@1082_d N_OUT6_Mp7@1082_g N_VDD_Mp7@1082_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1081 N_OUT7_Mn7@1081_d N_OUT6_Mn7@1081_g N_VSS_Mn7@1081_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1080 N_OUT7_Mn7@1080_d N_OUT6_Mn7@1080_g N_VSS_Mn7@1080_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1081 N_OUT7_Mp7@1081_d N_OUT6_Mp7@1081_g N_VDD_Mp7@1081_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1080 N_OUT7_Mp7@1080_d N_OUT6_Mp7@1080_g N_VDD_Mp7@1080_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1079 N_OUT7_Mn7@1079_d N_OUT6_Mn7@1079_g N_VSS_Mn7@1079_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1078 N_OUT7_Mn7@1078_d N_OUT6_Mn7@1078_g N_VSS_Mn7@1078_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1079 N_OUT7_Mp7@1079_d N_OUT6_Mp7@1079_g N_VDD_Mp7@1079_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1078 N_OUT7_Mp7@1078_d N_OUT6_Mp7@1078_g N_VDD_Mp7@1078_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1077 N_OUT7_Mn7@1077_d N_OUT6_Mn7@1077_g N_VSS_Mn7@1077_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1076 N_OUT7_Mn7@1076_d N_OUT6_Mn7@1076_g N_VSS_Mn7@1076_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1077 N_OUT7_Mp7@1077_d N_OUT6_Mp7@1077_g N_VDD_Mp7@1077_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1076 N_OUT7_Mp7@1076_d N_OUT6_Mp7@1076_g N_VDD_Mp7@1076_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1075 N_OUT7_Mn7@1075_d N_OUT6_Mn7@1075_g N_VSS_Mn7@1075_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1074 N_OUT7_Mn7@1074_d N_OUT6_Mn7@1074_g N_VSS_Mn7@1074_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1075 N_OUT7_Mp7@1075_d N_OUT6_Mp7@1075_g N_VDD_Mp7@1075_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1074 N_OUT7_Mp7@1074_d N_OUT6_Mp7@1074_g N_VDD_Mp7@1074_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1073 N_OUT7_Mn7@1073_d N_OUT6_Mn7@1073_g N_VSS_Mn7@1073_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1072 N_OUT7_Mn7@1072_d N_OUT6_Mn7@1072_g N_VSS_Mn7@1072_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1073 N_OUT7_Mp7@1073_d N_OUT6_Mp7@1073_g N_VDD_Mp7@1073_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1072 N_OUT7_Mp7@1072_d N_OUT6_Mp7@1072_g N_VDD_Mp7@1072_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1071 N_OUT7_Mn7@1071_d N_OUT6_Mn7@1071_g N_VSS_Mn7@1071_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1070 N_OUT7_Mn7@1070_d N_OUT6_Mn7@1070_g N_VSS_Mn7@1070_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1071 N_OUT7_Mp7@1071_d N_OUT6_Mp7@1071_g N_VDD_Mp7@1071_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1070 N_OUT7_Mp7@1070_d N_OUT6_Mp7@1070_g N_VDD_Mp7@1070_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1069 N_OUT7_Mn7@1069_d N_OUT6_Mn7@1069_g N_VSS_Mn7@1069_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1068 N_OUT7_Mn7@1068_d N_OUT6_Mn7@1068_g N_VSS_Mn7@1068_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1069 N_OUT7_Mp7@1069_d N_OUT6_Mp7@1069_g N_VDD_Mp7@1069_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1068 N_OUT7_Mp7@1068_d N_OUT6_Mp7@1068_g N_VDD_Mp7@1068_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1067 N_OUT7_Mn7@1067_d N_OUT6_Mn7@1067_g N_VSS_Mn7@1067_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1066 N_OUT7_Mn7@1066_d N_OUT6_Mn7@1066_g N_VSS_Mn7@1066_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1067 N_OUT7_Mp7@1067_d N_OUT6_Mp7@1067_g N_VDD_Mp7@1067_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1066 N_OUT7_Mp7@1066_d N_OUT6_Mp7@1066_g N_VDD_Mp7@1066_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1065 N_OUT7_Mn7@1065_d N_OUT6_Mn7@1065_g N_VSS_Mn7@1065_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1064 N_OUT7_Mn7@1064_d N_OUT6_Mn7@1064_g N_VSS_Mn7@1064_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1065 N_OUT7_Mp7@1065_d N_OUT6_Mp7@1065_g N_VDD_Mp7@1065_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1064 N_OUT7_Mp7@1064_d N_OUT6_Mp7@1064_g N_VDD_Mp7@1064_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1063 N_OUT7_Mn7@1063_d N_OUT6_Mn7@1063_g N_VSS_Mn7@1063_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1062 N_OUT7_Mn7@1062_d N_OUT6_Mn7@1062_g N_VSS_Mn7@1062_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1063 N_OUT7_Mp7@1063_d N_OUT6_Mp7@1063_g N_VDD_Mp7@1063_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1062 N_OUT7_Mp7@1062_d N_OUT6_Mp7@1062_g N_VDD_Mp7@1062_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1061 N_OUT7_Mn7@1061_d N_OUT6_Mn7@1061_g N_VSS_Mn7@1061_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1060 N_OUT7_Mn7@1060_d N_OUT6_Mn7@1060_g N_VSS_Mn7@1060_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1061 N_OUT7_Mp7@1061_d N_OUT6_Mp7@1061_g N_VDD_Mp7@1061_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1060 N_OUT7_Mp7@1060_d N_OUT6_Mp7@1060_g N_VDD_Mp7@1060_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1059 N_OUT7_Mn7@1059_d N_OUT6_Mn7@1059_g N_VSS_Mn7@1059_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1058 N_OUT7_Mn7@1058_d N_OUT6_Mn7@1058_g N_VSS_Mn7@1058_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1059 N_OUT7_Mp7@1059_d N_OUT6_Mp7@1059_g N_VDD_Mp7@1059_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1058 N_OUT7_Mp7@1058_d N_OUT6_Mp7@1058_g N_VDD_Mp7@1058_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1057 N_OUT7_Mn7@1057_d N_OUT6_Mn7@1057_g N_VSS_Mn7@1057_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1056 N_OUT7_Mn7@1056_d N_OUT6_Mn7@1056_g N_VSS_Mn7@1056_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1057 N_OUT7_Mp7@1057_d N_OUT6_Mp7@1057_g N_VDD_Mp7@1057_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1056 N_OUT7_Mp7@1056_d N_OUT6_Mp7@1056_g N_VDD_Mp7@1056_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1055 N_OUT7_Mn7@1055_d N_OUT6_Mn7@1055_g N_VSS_Mn7@1055_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1054 N_OUT7_Mn7@1054_d N_OUT6_Mn7@1054_g N_VSS_Mn7@1054_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1055 N_OUT7_Mp7@1055_d N_OUT6_Mp7@1055_g N_VDD_Mp7@1055_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1054 N_OUT7_Mp7@1054_d N_OUT6_Mp7@1054_g N_VDD_Mp7@1054_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1053 N_OUT7_Mn7@1053_d N_OUT6_Mn7@1053_g N_VSS_Mn7@1053_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1052 N_OUT7_Mn7@1052_d N_OUT6_Mn7@1052_g N_VSS_Mn7@1052_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1053 N_OUT7_Mp7@1053_d N_OUT6_Mp7@1053_g N_VDD_Mp7@1053_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1052 N_OUT7_Mp7@1052_d N_OUT6_Mp7@1052_g N_VDD_Mp7@1052_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1051 N_OUT7_Mn7@1051_d N_OUT6_Mn7@1051_g N_VSS_Mn7@1051_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1050 N_OUT7_Mn7@1050_d N_OUT6_Mn7@1050_g N_VSS_Mn7@1050_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1051 N_OUT7_Mp7@1051_d N_OUT6_Mp7@1051_g N_VDD_Mp7@1051_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1050 N_OUT7_Mp7@1050_d N_OUT6_Mp7@1050_g N_VDD_Mp7@1050_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1049 N_OUT7_Mn7@1049_d N_OUT6_Mn7@1049_g N_VSS_Mn7@1049_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1048 N_OUT7_Mn7@1048_d N_OUT6_Mn7@1048_g N_VSS_Mn7@1048_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1049 N_OUT7_Mp7@1049_d N_OUT6_Mp7@1049_g N_VDD_Mp7@1049_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1048 N_OUT7_Mp7@1048_d N_OUT6_Mp7@1048_g N_VDD_Mp7@1048_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1047 N_OUT7_Mn7@1047_d N_OUT6_Mn7@1047_g N_VSS_Mn7@1047_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1046 N_OUT7_Mn7@1046_d N_OUT6_Mn7@1046_g N_VSS_Mn7@1046_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1047 N_OUT7_Mp7@1047_d N_OUT6_Mp7@1047_g N_VDD_Mp7@1047_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1046 N_OUT7_Mp7@1046_d N_OUT6_Mp7@1046_g N_VDD_Mp7@1046_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1045 N_OUT7_Mn7@1045_d N_OUT6_Mn7@1045_g N_VSS_Mn7@1045_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1044 N_OUT7_Mn7@1044_d N_OUT6_Mn7@1044_g N_VSS_Mn7@1044_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1045 N_OUT7_Mp7@1045_d N_OUT6_Mp7@1045_g N_VDD_Mp7@1045_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1044 N_OUT7_Mp7@1044_d N_OUT6_Mp7@1044_g N_VDD_Mp7@1044_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1043 N_OUT7_Mn7@1043_d N_OUT6_Mn7@1043_g N_VSS_Mn7@1043_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1042 N_OUT7_Mn7@1042_d N_OUT6_Mn7@1042_g N_VSS_Mn7@1042_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1043 N_OUT7_Mp7@1043_d N_OUT6_Mp7@1043_g N_VDD_Mp7@1043_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1042 N_OUT7_Mp7@1042_d N_OUT6_Mp7@1042_g N_VDD_Mp7@1042_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1041 N_OUT7_Mn7@1041_d N_OUT6_Mn7@1041_g N_VSS_Mn7@1041_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1040 N_OUT7_Mn7@1040_d N_OUT6_Mn7@1040_g N_VSS_Mn7@1040_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1041 N_OUT7_Mp7@1041_d N_OUT6_Mp7@1041_g N_VDD_Mp7@1041_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1040 N_OUT7_Mp7@1040_d N_OUT6_Mp7@1040_g N_VDD_Mp7@1040_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1039 N_OUT7_Mn7@1039_d N_OUT6_Mn7@1039_g N_VSS_Mn7@1039_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1038 N_OUT7_Mn7@1038_d N_OUT6_Mn7@1038_g N_VSS_Mn7@1038_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1039 N_OUT7_Mp7@1039_d N_OUT6_Mp7@1039_g N_VDD_Mp7@1039_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1038 N_OUT7_Mp7@1038_d N_OUT6_Mp7@1038_g N_VDD_Mp7@1038_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1037 N_OUT7_Mn7@1037_d N_OUT6_Mn7@1037_g N_VSS_Mn7@1037_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1036 N_OUT7_Mn7@1036_d N_OUT6_Mn7@1036_g N_VSS_Mn7@1036_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1037 N_OUT7_Mp7@1037_d N_OUT6_Mp7@1037_g N_VDD_Mp7@1037_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1036 N_OUT7_Mp7@1036_d N_OUT6_Mp7@1036_g N_VDD_Mp7@1036_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1035 N_OUT7_Mn7@1035_d N_OUT6_Mn7@1035_g N_VSS_Mn7@1035_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1034 N_OUT7_Mn7@1034_d N_OUT6_Mn7@1034_g N_VSS_Mn7@1034_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1035 N_OUT7_Mp7@1035_d N_OUT6_Mp7@1035_g N_VDD_Mp7@1035_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1034 N_OUT7_Mp7@1034_d N_OUT6_Mp7@1034_g N_VDD_Mp7@1034_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1033 N_OUT7_Mn7@1033_d N_OUT6_Mn7@1033_g N_VSS_Mn7@1033_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1032 N_OUT7_Mn7@1032_d N_OUT6_Mn7@1032_g N_VSS_Mn7@1032_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1033 N_OUT7_Mp7@1033_d N_OUT6_Mp7@1033_g N_VDD_Mp7@1033_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1032 N_OUT7_Mp7@1032_d N_OUT6_Mp7@1032_g N_VDD_Mp7@1032_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1031 N_OUT7_Mn7@1031_d N_OUT6_Mn7@1031_g N_VSS_Mn7@1031_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1030 N_OUT7_Mn7@1030_d N_OUT6_Mn7@1030_g N_VSS_Mn7@1030_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1031 N_OUT7_Mp7@1031_d N_OUT6_Mp7@1031_g N_VDD_Mp7@1031_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1030 N_OUT7_Mp7@1030_d N_OUT6_Mp7@1030_g N_VDD_Mp7@1030_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1029 N_OUT7_Mn7@1029_d N_OUT6_Mn7@1029_g N_VSS_Mn7@1029_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1028 N_OUT7_Mn7@1028_d N_OUT6_Mn7@1028_g N_VSS_Mn7@1028_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1029 N_OUT7_Mp7@1029_d N_OUT6_Mp7@1029_g N_VDD_Mp7@1029_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1028 N_OUT7_Mp7@1028_d N_OUT6_Mp7@1028_g N_VDD_Mp7@1028_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1027 N_OUT7_Mn7@1027_d N_OUT6_Mn7@1027_g N_VSS_Mn7@1027_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1026 N_OUT7_Mn7@1026_d N_OUT6_Mn7@1026_g N_VSS_Mn7@1026_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1027 N_OUT7_Mp7@1027_d N_OUT6_Mp7@1027_g N_VDD_Mp7@1027_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1026 N_OUT7_Mp7@1026_d N_OUT6_Mp7@1026_g N_VDD_Mp7@1026_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3713 N_OUT8_Mn8@3713_d N_OUT7_Mn8@3713_g N_VSS_Mn8@3713_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3712 N_OUT8_Mn8@3712_d N_OUT7_Mn8@3712_g N_VSS_Mn8@3712_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3713 N_OUT8_Mp8@3713_d N_OUT7_Mp8@3713_g N_VDD_Mp8@3713_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3712 N_OUT8_Mp8@3712_d N_OUT7_Mp8@3712_g N_VDD_Mp8@3712_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3711 N_OUT8_Mn8@3711_d N_OUT7_Mn8@3711_g N_VSS_Mn8@3711_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3710 N_OUT8_Mn8@3710_d N_OUT7_Mn8@3710_g N_VSS_Mn8@3710_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3711 N_OUT8_Mp8@3711_d N_OUT7_Mp8@3711_g N_VDD_Mp8@3711_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3710 N_OUT8_Mp8@3710_d N_OUT7_Mp8@3710_g N_VDD_Mp8@3710_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3709 N_OUT8_Mn8@3709_d N_OUT7_Mn8@3709_g N_VSS_Mn8@3709_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3708 N_OUT8_Mn8@3708_d N_OUT7_Mn8@3708_g N_VSS_Mn8@3708_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3709 N_OUT8_Mp8@3709_d N_OUT7_Mp8@3709_g N_VDD_Mp8@3709_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3708 N_OUT8_Mp8@3708_d N_OUT7_Mp8@3708_g N_VDD_Mp8@3708_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3707 N_OUT8_Mn8@3707_d N_OUT7_Mn8@3707_g N_VSS_Mn8@3707_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3706 N_OUT8_Mn8@3706_d N_OUT7_Mn8@3706_g N_VSS_Mn8@3706_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3707 N_OUT8_Mp8@3707_d N_OUT7_Mp8@3707_g N_VDD_Mp8@3707_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3706 N_OUT8_Mp8@3706_d N_OUT7_Mp8@3706_g N_VDD_Mp8@3706_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3705 N_OUT8_Mn8@3705_d N_OUT7_Mn8@3705_g N_VSS_Mn8@3705_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3704 N_OUT8_Mn8@3704_d N_OUT7_Mn8@3704_g N_VSS_Mn8@3704_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3705 N_OUT8_Mp8@3705_d N_OUT7_Mp8@3705_g N_VDD_Mp8@3705_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3704 N_OUT8_Mp8@3704_d N_OUT7_Mp8@3704_g N_VDD_Mp8@3704_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3703 N_OUT8_Mn8@3703_d N_OUT7_Mn8@3703_g N_VSS_Mn8@3703_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3702 N_OUT8_Mn8@3702_d N_OUT7_Mn8@3702_g N_VSS_Mn8@3702_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3703 N_OUT8_Mp8@3703_d N_OUT7_Mp8@3703_g N_VDD_Mp8@3703_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3702 N_OUT8_Mp8@3702_d N_OUT7_Mp8@3702_g N_VDD_Mp8@3702_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3701 N_OUT8_Mn8@3701_d N_OUT7_Mn8@3701_g N_VSS_Mn8@3701_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3700 N_OUT8_Mn8@3700_d N_OUT7_Mn8@3700_g N_VSS_Mn8@3700_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3701 N_OUT8_Mp8@3701_d N_OUT7_Mp8@3701_g N_VDD_Mp8@3701_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3700 N_OUT8_Mp8@3700_d N_OUT7_Mp8@3700_g N_VDD_Mp8@3700_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3699 N_OUT8_Mn8@3699_d N_OUT7_Mn8@3699_g N_VSS_Mn8@3699_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3698 N_OUT8_Mn8@3698_d N_OUT7_Mn8@3698_g N_VSS_Mn8@3698_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3699 N_OUT8_Mp8@3699_d N_OUT7_Mp8@3699_g N_VDD_Mp8@3699_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3698 N_OUT8_Mp8@3698_d N_OUT7_Mp8@3698_g N_VDD_Mp8@3698_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3697 N_OUT8_Mn8@3697_d N_OUT7_Mn8@3697_g N_VSS_Mn8@3697_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3696 N_OUT8_Mn8@3696_d N_OUT7_Mn8@3696_g N_VSS_Mn8@3696_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3697 N_OUT8_Mp8@3697_d N_OUT7_Mp8@3697_g N_VDD_Mp8@3697_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3696 N_OUT8_Mp8@3696_d N_OUT7_Mp8@3696_g N_VDD_Mp8@3696_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3695 N_OUT8_Mn8@3695_d N_OUT7_Mn8@3695_g N_VSS_Mn8@3695_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3694 N_OUT8_Mn8@3694_d N_OUT7_Mn8@3694_g N_VSS_Mn8@3694_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3695 N_OUT8_Mp8@3695_d N_OUT7_Mp8@3695_g N_VDD_Mp8@3695_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3694 N_OUT8_Mp8@3694_d N_OUT7_Mp8@3694_g N_VDD_Mp8@3694_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3693 N_OUT8_Mn8@3693_d N_OUT7_Mn8@3693_g N_VSS_Mn8@3693_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3692 N_OUT8_Mn8@3692_d N_OUT7_Mn8@3692_g N_VSS_Mn8@3692_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3693 N_OUT8_Mp8@3693_d N_OUT7_Mp8@3693_g N_VDD_Mp8@3693_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3692 N_OUT8_Mp8@3692_d N_OUT7_Mp8@3692_g N_VDD_Mp8@3692_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3691 N_OUT8_Mn8@3691_d N_OUT7_Mn8@3691_g N_VSS_Mn8@3691_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3690 N_OUT8_Mn8@3690_d N_OUT7_Mn8@3690_g N_VSS_Mn8@3690_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3691 N_OUT8_Mp8@3691_d N_OUT7_Mp8@3691_g N_VDD_Mp8@3691_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3690 N_OUT8_Mp8@3690_d N_OUT7_Mp8@3690_g N_VDD_Mp8@3690_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3689 N_OUT8_Mn8@3689_d N_OUT7_Mn8@3689_g N_VSS_Mn8@3689_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3688 N_OUT8_Mn8@3688_d N_OUT7_Mn8@3688_g N_VSS_Mn8@3688_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3689 N_OUT8_Mp8@3689_d N_OUT7_Mp8@3689_g N_VDD_Mp8@3689_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3688 N_OUT8_Mp8@3688_d N_OUT7_Mp8@3688_g N_VDD_Mp8@3688_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3687 N_OUT8_Mn8@3687_d N_OUT7_Mn8@3687_g N_VSS_Mn8@3687_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3686 N_OUT8_Mn8@3686_d N_OUT7_Mn8@3686_g N_VSS_Mn8@3686_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3687 N_OUT8_Mp8@3687_d N_OUT7_Mp8@3687_g N_VDD_Mp8@3687_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3686 N_OUT8_Mp8@3686_d N_OUT7_Mp8@3686_g N_VDD_Mp8@3686_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3685 N_OUT8_Mn8@3685_d N_OUT7_Mn8@3685_g N_VSS_Mn8@3685_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3684 N_OUT8_Mn8@3684_d N_OUT7_Mn8@3684_g N_VSS_Mn8@3684_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3685 N_OUT8_Mp8@3685_d N_OUT7_Mp8@3685_g N_VDD_Mp8@3685_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3684 N_OUT8_Mp8@3684_d N_OUT7_Mp8@3684_g N_VDD_Mp8@3684_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3683 N_OUT8_Mn8@3683_d N_OUT7_Mn8@3683_g N_VSS_Mn8@3683_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3682 N_OUT8_Mn8@3682_d N_OUT7_Mn8@3682_g N_VSS_Mn8@3682_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3683 N_OUT8_Mp8@3683_d N_OUT7_Mp8@3683_g N_VDD_Mp8@3683_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3682 N_OUT8_Mp8@3682_d N_OUT7_Mp8@3682_g N_VDD_Mp8@3682_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3681 N_OUT8_Mn8@3681_d N_OUT7_Mn8@3681_g N_VSS_Mn8@3681_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3680 N_OUT8_Mn8@3680_d N_OUT7_Mn8@3680_g N_VSS_Mn8@3680_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3681 N_OUT8_Mp8@3681_d N_OUT7_Mp8@3681_g N_VDD_Mp8@3681_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3680 N_OUT8_Mp8@3680_d N_OUT7_Mp8@3680_g N_VDD_Mp8@3680_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3679 N_OUT8_Mn8@3679_d N_OUT7_Mn8@3679_g N_VSS_Mn8@3679_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3678 N_OUT8_Mn8@3678_d N_OUT7_Mn8@3678_g N_VSS_Mn8@3678_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3679 N_OUT8_Mp8@3679_d N_OUT7_Mp8@3679_g N_VDD_Mp8@3679_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3678 N_OUT8_Mp8@3678_d N_OUT7_Mp8@3678_g N_VDD_Mp8@3678_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3677 N_OUT8_Mn8@3677_d N_OUT7_Mn8@3677_g N_VSS_Mn8@3677_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3676 N_OUT8_Mn8@3676_d N_OUT7_Mn8@3676_g N_VSS_Mn8@3676_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3677 N_OUT8_Mp8@3677_d N_OUT7_Mp8@3677_g N_VDD_Mp8@3677_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3676 N_OUT8_Mp8@3676_d N_OUT7_Mp8@3676_g N_VDD_Mp8@3676_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3675 N_OUT8_Mn8@3675_d N_OUT7_Mn8@3675_g N_VSS_Mn8@3675_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3674 N_OUT8_Mn8@3674_d N_OUT7_Mn8@3674_g N_VSS_Mn8@3674_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3675 N_OUT8_Mp8@3675_d N_OUT7_Mp8@3675_g N_VDD_Mp8@3675_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3674 N_OUT8_Mp8@3674_d N_OUT7_Mp8@3674_g N_VDD_Mp8@3674_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3673 N_OUT8_Mn8@3673_d N_OUT7_Mn8@3673_g N_VSS_Mn8@3673_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3672 N_OUT8_Mn8@3672_d N_OUT7_Mn8@3672_g N_VSS_Mn8@3672_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3673 N_OUT8_Mp8@3673_d N_OUT7_Mp8@3673_g N_VDD_Mp8@3673_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3672 N_OUT8_Mp8@3672_d N_OUT7_Mp8@3672_g N_VDD_Mp8@3672_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3671 N_OUT8_Mn8@3671_d N_OUT7_Mn8@3671_g N_VSS_Mn8@3671_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3670 N_OUT8_Mn8@3670_d N_OUT7_Mn8@3670_g N_VSS_Mn8@3670_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3671 N_OUT8_Mp8@3671_d N_OUT7_Mp8@3671_g N_VDD_Mp8@3671_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3670 N_OUT8_Mp8@3670_d N_OUT7_Mp8@3670_g N_VDD_Mp8@3670_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3669 N_OUT8_Mn8@3669_d N_OUT7_Mn8@3669_g N_VSS_Mn8@3669_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3668 N_OUT8_Mn8@3668_d N_OUT7_Mn8@3668_g N_VSS_Mn8@3668_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3669 N_OUT8_Mp8@3669_d N_OUT7_Mp8@3669_g N_VDD_Mp8@3669_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3668 N_OUT8_Mp8@3668_d N_OUT7_Mp8@3668_g N_VDD_Mp8@3668_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3667 N_OUT8_Mn8@3667_d N_OUT7_Mn8@3667_g N_VSS_Mn8@3667_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3666 N_OUT8_Mn8@3666_d N_OUT7_Mn8@3666_g N_VSS_Mn8@3666_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3667 N_OUT8_Mp8@3667_d N_OUT7_Mp8@3667_g N_VDD_Mp8@3667_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3666 N_OUT8_Mp8@3666_d N_OUT7_Mp8@3666_g N_VDD_Mp8@3666_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3665 N_OUT8_Mn8@3665_d N_OUT7_Mn8@3665_g N_VSS_Mn8@3665_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3664 N_OUT8_Mn8@3664_d N_OUT7_Mn8@3664_g N_VSS_Mn8@3664_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3665 N_OUT8_Mp8@3665_d N_OUT7_Mp8@3665_g N_VDD_Mp8@3665_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3664 N_OUT8_Mp8@3664_d N_OUT7_Mp8@3664_g N_VDD_Mp8@3664_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3663 N_OUT8_Mn8@3663_d N_OUT7_Mn8@3663_g N_VSS_Mn8@3663_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3662 N_OUT8_Mn8@3662_d N_OUT7_Mn8@3662_g N_VSS_Mn8@3662_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3663 N_OUT8_Mp8@3663_d N_OUT7_Mp8@3663_g N_VDD_Mp8@3663_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3662 N_OUT8_Mp8@3662_d N_OUT7_Mp8@3662_g N_VDD_Mp8@3662_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3661 N_OUT8_Mn8@3661_d N_OUT7_Mn8@3661_g N_VSS_Mn8@3661_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3660 N_OUT8_Mn8@3660_d N_OUT7_Mn8@3660_g N_VSS_Mn8@3660_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3661 N_OUT8_Mp8@3661_d N_OUT7_Mp8@3661_g N_VDD_Mp8@3661_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3660 N_OUT8_Mp8@3660_d N_OUT7_Mp8@3660_g N_VDD_Mp8@3660_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3659 N_OUT8_Mn8@3659_d N_OUT7_Mn8@3659_g N_VSS_Mn8@3659_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3658 N_OUT8_Mn8@3658_d N_OUT7_Mn8@3658_g N_VSS_Mn8@3658_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3659 N_OUT8_Mp8@3659_d N_OUT7_Mp8@3659_g N_VDD_Mp8@3659_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3658 N_OUT8_Mp8@3658_d N_OUT7_Mp8@3658_g N_VDD_Mp8@3658_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3657 N_OUT8_Mn8@3657_d N_OUT7_Mn8@3657_g N_VSS_Mn8@3657_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3656 N_OUT8_Mn8@3656_d N_OUT7_Mn8@3656_g N_VSS_Mn8@3656_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3657 N_OUT8_Mp8@3657_d N_OUT7_Mp8@3657_g N_VDD_Mp8@3657_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3656 N_OUT8_Mp8@3656_d N_OUT7_Mp8@3656_g N_VDD_Mp8@3656_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3655 N_OUT8_Mn8@3655_d N_OUT7_Mn8@3655_g N_VSS_Mn8@3655_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3654 N_OUT8_Mn8@3654_d N_OUT7_Mn8@3654_g N_VSS_Mn8@3654_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3655 N_OUT8_Mp8@3655_d N_OUT7_Mp8@3655_g N_VDD_Mp8@3655_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3654 N_OUT8_Mp8@3654_d N_OUT7_Mp8@3654_g N_VDD_Mp8@3654_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3653 N_OUT8_Mn8@3653_d N_OUT7_Mn8@3653_g N_VSS_Mn8@3653_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3652 N_OUT8_Mn8@3652_d N_OUT7_Mn8@3652_g N_VSS_Mn8@3652_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3653 N_OUT8_Mp8@3653_d N_OUT7_Mp8@3653_g N_VDD_Mp8@3653_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3652 N_OUT8_Mp8@3652_d N_OUT7_Mp8@3652_g N_VDD_Mp8@3652_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3651 N_OUT8_Mn8@3651_d N_OUT7_Mn8@3651_g N_VSS_Mn8@3651_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3650 N_OUT8_Mn8@3650_d N_OUT7_Mn8@3650_g N_VSS_Mn8@3650_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3651 N_OUT8_Mp8@3651_d N_OUT7_Mp8@3651_g N_VDD_Mp8@3651_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3650 N_OUT8_Mp8@3650_d N_OUT7_Mp8@3650_g N_VDD_Mp8@3650_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3649 N_OUT8_Mn8@3649_d N_OUT7_Mn8@3649_g N_VSS_Mn8@3649_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3648 N_OUT8_Mn8@3648_d N_OUT7_Mn8@3648_g N_VSS_Mn8@3648_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3649 N_OUT8_Mp8@3649_d N_OUT7_Mp8@3649_g N_VDD_Mp8@3649_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3648 N_OUT8_Mp8@3648_d N_OUT7_Mp8@3648_g N_VDD_Mp8@3648_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3647 N_OUT8_Mn8@3647_d N_OUT7_Mn8@3647_g N_VSS_Mn8@3647_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3646 N_OUT8_Mn8@3646_d N_OUT7_Mn8@3646_g N_VSS_Mn8@3646_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3647 N_OUT8_Mp8@3647_d N_OUT7_Mp8@3647_g N_VDD_Mp8@3647_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3646 N_OUT8_Mp8@3646_d N_OUT7_Mp8@3646_g N_VDD_Mp8@3646_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3645 N_OUT8_Mn8@3645_d N_OUT7_Mn8@3645_g N_VSS_Mn8@3645_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3644 N_OUT8_Mn8@3644_d N_OUT7_Mn8@3644_g N_VSS_Mn8@3644_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3645 N_OUT8_Mp8@3645_d N_OUT7_Mp8@3645_g N_VDD_Mp8@3645_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3644 N_OUT8_Mp8@3644_d N_OUT7_Mp8@3644_g N_VDD_Mp8@3644_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3643 N_OUT8_Mn8@3643_d N_OUT7_Mn8@3643_g N_VSS_Mn8@3643_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3642 N_OUT8_Mn8@3642_d N_OUT7_Mn8@3642_g N_VSS_Mn8@3642_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3643 N_OUT8_Mp8@3643_d N_OUT7_Mp8@3643_g N_VDD_Mp8@3643_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3642 N_OUT8_Mp8@3642_d N_OUT7_Mp8@3642_g N_VDD_Mp8@3642_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3641 N_OUT8_Mn8@3641_d N_OUT7_Mn8@3641_g N_VSS_Mn8@3641_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3640 N_OUT8_Mn8@3640_d N_OUT7_Mn8@3640_g N_VSS_Mn8@3640_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3641 N_OUT8_Mp8@3641_d N_OUT7_Mp8@3641_g N_VDD_Mp8@3641_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3640 N_OUT8_Mp8@3640_d N_OUT7_Mp8@3640_g N_VDD_Mp8@3640_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3639 N_OUT8_Mn8@3639_d N_OUT7_Mn8@3639_g N_VSS_Mn8@3639_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3638 N_OUT8_Mn8@3638_d N_OUT7_Mn8@3638_g N_VSS_Mn8@3638_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3639 N_OUT8_Mp8@3639_d N_OUT7_Mp8@3639_g N_VDD_Mp8@3639_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3638 N_OUT8_Mp8@3638_d N_OUT7_Mp8@3638_g N_VDD_Mp8@3638_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3637 N_OUT8_Mn8@3637_d N_OUT7_Mn8@3637_g N_VSS_Mn8@3637_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3636 N_OUT8_Mn8@3636_d N_OUT7_Mn8@3636_g N_VSS_Mn8@3636_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3637 N_OUT8_Mp8@3637_d N_OUT7_Mp8@3637_g N_VDD_Mp8@3637_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3636 N_OUT8_Mp8@3636_d N_OUT7_Mp8@3636_g N_VDD_Mp8@3636_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3635 N_OUT8_Mn8@3635_d N_OUT7_Mn8@3635_g N_VSS_Mn8@3635_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3634 N_OUT8_Mn8@3634_d N_OUT7_Mn8@3634_g N_VSS_Mn8@3634_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3635 N_OUT8_Mp8@3635_d N_OUT7_Mp8@3635_g N_VDD_Mp8@3635_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3634 N_OUT8_Mp8@3634_d N_OUT7_Mp8@3634_g N_VDD_Mp8@3634_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3633 N_OUT8_Mn8@3633_d N_OUT7_Mn8@3633_g N_VSS_Mn8@3633_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3632 N_OUT8_Mn8@3632_d N_OUT7_Mn8@3632_g N_VSS_Mn8@3632_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3633 N_OUT8_Mp8@3633_d N_OUT7_Mp8@3633_g N_VDD_Mp8@3633_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3632 N_OUT8_Mp8@3632_d N_OUT7_Mp8@3632_g N_VDD_Mp8@3632_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3631 N_OUT8_Mn8@3631_d N_OUT7_Mn8@3631_g N_VSS_Mn8@3631_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3630 N_OUT8_Mn8@3630_d N_OUT7_Mn8@3630_g N_VSS_Mn8@3630_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3631 N_OUT8_Mp8@3631_d N_OUT7_Mp8@3631_g N_VDD_Mp8@3631_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3630 N_OUT8_Mp8@3630_d N_OUT7_Mp8@3630_g N_VDD_Mp8@3630_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3629 N_OUT8_Mn8@3629_d N_OUT7_Mn8@3629_g N_VSS_Mn8@3629_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3628 N_OUT8_Mn8@3628_d N_OUT7_Mn8@3628_g N_VSS_Mn8@3628_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3629 N_OUT8_Mp8@3629_d N_OUT7_Mp8@3629_g N_VDD_Mp8@3629_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3628 N_OUT8_Mp8@3628_d N_OUT7_Mp8@3628_g N_VDD_Mp8@3628_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3627 N_OUT8_Mn8@3627_d N_OUT7_Mn8@3627_g N_VSS_Mn8@3627_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3626 N_OUT8_Mn8@3626_d N_OUT7_Mn8@3626_g N_VSS_Mn8@3626_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3627 N_OUT8_Mp8@3627_d N_OUT7_Mp8@3627_g N_VDD_Mp8@3627_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3626 N_OUT8_Mp8@3626_d N_OUT7_Mp8@3626_g N_VDD_Mp8@3626_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3625 N_OUT8_Mn8@3625_d N_OUT7_Mn8@3625_g N_VSS_Mn8@3625_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3624 N_OUT8_Mn8@3624_d N_OUT7_Mn8@3624_g N_VSS_Mn8@3624_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3625 N_OUT8_Mp8@3625_d N_OUT7_Mp8@3625_g N_VDD_Mp8@3625_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3624 N_OUT8_Mp8@3624_d N_OUT7_Mp8@3624_g N_VDD_Mp8@3624_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3623 N_OUT8_Mn8@3623_d N_OUT7_Mn8@3623_g N_VSS_Mn8@3623_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3622 N_OUT8_Mn8@3622_d N_OUT7_Mn8@3622_g N_VSS_Mn8@3622_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3623 N_OUT8_Mp8@3623_d N_OUT7_Mp8@3623_g N_VDD_Mp8@3623_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3622 N_OUT8_Mp8@3622_d N_OUT7_Mp8@3622_g N_VDD_Mp8@3622_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3621 N_OUT8_Mn8@3621_d N_OUT7_Mn8@3621_g N_VSS_Mn8@3621_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3620 N_OUT8_Mn8@3620_d N_OUT7_Mn8@3620_g N_VSS_Mn8@3620_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3621 N_OUT8_Mp8@3621_d N_OUT7_Mp8@3621_g N_VDD_Mp8@3621_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3620 N_OUT8_Mp8@3620_d N_OUT7_Mp8@3620_g N_VDD_Mp8@3620_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3619 N_OUT8_Mn8@3619_d N_OUT7_Mn8@3619_g N_VSS_Mn8@3619_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3618 N_OUT8_Mn8@3618_d N_OUT7_Mn8@3618_g N_VSS_Mn8@3618_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3619 N_OUT8_Mp8@3619_d N_OUT7_Mp8@3619_g N_VDD_Mp8@3619_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3618 N_OUT8_Mp8@3618_d N_OUT7_Mp8@3618_g N_VDD_Mp8@3618_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3617 N_OUT8_Mn8@3617_d N_OUT7_Mn8@3617_g N_VSS_Mn8@3617_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3616 N_OUT8_Mn8@3616_d N_OUT7_Mn8@3616_g N_VSS_Mn8@3616_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3617 N_OUT8_Mp8@3617_d N_OUT7_Mp8@3617_g N_VDD_Mp8@3617_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3616 N_OUT8_Mp8@3616_d N_OUT7_Mp8@3616_g N_VDD_Mp8@3616_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3615 N_OUT8_Mn8@3615_d N_OUT7_Mn8@3615_g N_VSS_Mn8@3615_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3614 N_OUT8_Mn8@3614_d N_OUT7_Mn8@3614_g N_VSS_Mn8@3614_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3615 N_OUT8_Mp8@3615_d N_OUT7_Mp8@3615_g N_VDD_Mp8@3615_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3614 N_OUT8_Mp8@3614_d N_OUT7_Mp8@3614_g N_VDD_Mp8@3614_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3613 N_OUT8_Mn8@3613_d N_OUT7_Mn8@3613_g N_VSS_Mn8@3613_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3612 N_OUT8_Mn8@3612_d N_OUT7_Mn8@3612_g N_VSS_Mn8@3612_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3613 N_OUT8_Mp8@3613_d N_OUT7_Mp8@3613_g N_VDD_Mp8@3613_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3612 N_OUT8_Mp8@3612_d N_OUT7_Mp8@3612_g N_VDD_Mp8@3612_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3611 N_OUT8_Mn8@3611_d N_OUT7_Mn8@3611_g N_VSS_Mn8@3611_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3610 N_OUT8_Mn8@3610_d N_OUT7_Mn8@3610_g N_VSS_Mn8@3610_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3611 N_OUT8_Mp8@3611_d N_OUT7_Mp8@3611_g N_VDD_Mp8@3611_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3610 N_OUT8_Mp8@3610_d N_OUT7_Mp8@3610_g N_VDD_Mp8@3610_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3609 N_OUT8_Mn8@3609_d N_OUT7_Mn8@3609_g N_VSS_Mn8@3609_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3608 N_OUT8_Mn8@3608_d N_OUT7_Mn8@3608_g N_VSS_Mn8@3608_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3609 N_OUT8_Mp8@3609_d N_OUT7_Mp8@3609_g N_VDD_Mp8@3609_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3608 N_OUT8_Mp8@3608_d N_OUT7_Mp8@3608_g N_VDD_Mp8@3608_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3607 N_OUT8_Mn8@3607_d N_OUT7_Mn8@3607_g N_VSS_Mn8@3607_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3606 N_OUT8_Mn8@3606_d N_OUT7_Mn8@3606_g N_VSS_Mn8@3606_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3607 N_OUT8_Mp8@3607_d N_OUT7_Mp8@3607_g N_VDD_Mp8@3607_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3606 N_OUT8_Mp8@3606_d N_OUT7_Mp8@3606_g N_VDD_Mp8@3606_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3605 N_OUT8_Mn8@3605_d N_OUT7_Mn8@3605_g N_VSS_Mn8@3605_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3604 N_OUT8_Mn8@3604_d N_OUT7_Mn8@3604_g N_VSS_Mn8@3604_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3605 N_OUT8_Mp8@3605_d N_OUT7_Mp8@3605_g N_VDD_Mp8@3605_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3604 N_OUT8_Mp8@3604_d N_OUT7_Mp8@3604_g N_VDD_Mp8@3604_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3603 N_OUT8_Mn8@3603_d N_OUT7_Mn8@3603_g N_VSS_Mn8@3603_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3602 N_OUT8_Mn8@3602_d N_OUT7_Mn8@3602_g N_VSS_Mn8@3602_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3603 N_OUT8_Mp8@3603_d N_OUT7_Mp8@3603_g N_VDD_Mp8@3603_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3602 N_OUT8_Mp8@3602_d N_OUT7_Mp8@3602_g N_VDD_Mp8@3602_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3601 N_OUT8_Mn8@3601_d N_OUT7_Mn8@3601_g N_VSS_Mn8@3601_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3600 N_OUT8_Mn8@3600_d N_OUT7_Mn8@3600_g N_VSS_Mn8@3600_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3601 N_OUT8_Mp8@3601_d N_OUT7_Mp8@3601_g N_VDD_Mp8@3601_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3600 N_OUT8_Mp8@3600_d N_OUT7_Mp8@3600_g N_VDD_Mp8@3600_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3599 N_OUT8_Mn8@3599_d N_OUT7_Mn8@3599_g N_VSS_Mn8@3599_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3598 N_OUT8_Mn8@3598_d N_OUT7_Mn8@3598_g N_VSS_Mn8@3598_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3599 N_OUT8_Mp8@3599_d N_OUT7_Mp8@3599_g N_VDD_Mp8@3599_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3598 N_OUT8_Mp8@3598_d N_OUT7_Mp8@3598_g N_VDD_Mp8@3598_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3597 N_OUT8_Mn8@3597_d N_OUT7_Mn8@3597_g N_VSS_Mn8@3597_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3596 N_OUT8_Mn8@3596_d N_OUT7_Mn8@3596_g N_VSS_Mn8@3596_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3597 N_OUT8_Mp8@3597_d N_OUT7_Mp8@3597_g N_VDD_Mp8@3597_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3596 N_OUT8_Mp8@3596_d N_OUT7_Mp8@3596_g N_VDD_Mp8@3596_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3595 N_OUT8_Mn8@3595_d N_OUT7_Mn8@3595_g N_VSS_Mn8@3595_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3594 N_OUT8_Mn8@3594_d N_OUT7_Mn8@3594_g N_VSS_Mn8@3594_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3595 N_OUT8_Mp8@3595_d N_OUT7_Mp8@3595_g N_VDD_Mp8@3595_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3594 N_OUT8_Mp8@3594_d N_OUT7_Mp8@3594_g N_VDD_Mp8@3594_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3593 N_OUT8_Mn8@3593_d N_OUT7_Mn8@3593_g N_VSS_Mn8@3593_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3592 N_OUT8_Mn8@3592_d N_OUT7_Mn8@3592_g N_VSS_Mn8@3592_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3593 N_OUT8_Mp8@3593_d N_OUT7_Mp8@3593_g N_VDD_Mp8@3593_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3592 N_OUT8_Mp8@3592_d N_OUT7_Mp8@3592_g N_VDD_Mp8@3592_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3591 N_OUT8_Mn8@3591_d N_OUT7_Mn8@3591_g N_VSS_Mn8@3591_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3590 N_OUT8_Mn8@3590_d N_OUT7_Mn8@3590_g N_VSS_Mn8@3590_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3591 N_OUT8_Mp8@3591_d N_OUT7_Mp8@3591_g N_VDD_Mp8@3591_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3590 N_OUT8_Mp8@3590_d N_OUT7_Mp8@3590_g N_VDD_Mp8@3590_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3589 N_OUT8_Mn8@3589_d N_OUT7_Mn8@3589_g N_VSS_Mn8@3589_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3588 N_OUT8_Mn8@3588_d N_OUT7_Mn8@3588_g N_VSS_Mn8@3588_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3589 N_OUT8_Mp8@3589_d N_OUT7_Mp8@3589_g N_VDD_Mp8@3589_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3588 N_OUT8_Mp8@3588_d N_OUT7_Mp8@3588_g N_VDD_Mp8@3588_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3587 N_OUT8_Mn8@3587_d N_OUT7_Mn8@3587_g N_VSS_Mn8@3587_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3586 N_OUT8_Mn8@3586_d N_OUT7_Mn8@3586_g N_VSS_Mn8@3586_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3587 N_OUT8_Mp8@3587_d N_OUT7_Mp8@3587_g N_VDD_Mp8@3587_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3586 N_OUT8_Mp8@3586_d N_OUT7_Mp8@3586_g N_VDD_Mp8@3586_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4995 N_OUT9_Mn9@4995_d N_OUT8_Mn9@4995_g N_VSS_Mn9@4995_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4994 N_OUT9_Mn9@4994_d N_OUT8_Mn9@4994_g N_VSS_Mn9@4994_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4995 N_OUT9_Mp9@4995_d N_OUT8_Mp9@4995_g N_VDD_Mp9@4995_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4994 N_OUT9_Mp9@4994_d N_OUT8_Mp9@4994_g N_VDD_Mp9@4994_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4993 N_OUT9_Mn9@4993_d N_OUT8_Mn9@4993_g N_VSS_Mn9@4993_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4992 N_OUT9_Mn9@4992_d N_OUT8_Mn9@4992_g N_VSS_Mn9@4992_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4993 N_OUT9_Mp9@4993_d N_OUT8_Mp9@4993_g N_VDD_Mp9@4993_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4992 N_OUT9_Mp9@4992_d N_OUT8_Mp9@4992_g N_VDD_Mp9@4992_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4991 N_OUT9_Mn9@4991_d N_OUT8_Mn9@4991_g N_VSS_Mn9@4991_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4990 N_OUT9_Mn9@4990_d N_OUT8_Mn9@4990_g N_VSS_Mn9@4990_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4991 N_OUT9_Mp9@4991_d N_OUT8_Mp9@4991_g N_VDD_Mp9@4991_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4990 N_OUT9_Mp9@4990_d N_OUT8_Mp9@4990_g N_VDD_Mp9@4990_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4989 N_OUT9_Mn9@4989_d N_OUT8_Mn9@4989_g N_VSS_Mn9@4989_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4988 N_OUT9_Mn9@4988_d N_OUT8_Mn9@4988_g N_VSS_Mn9@4988_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4989 N_OUT9_Mp9@4989_d N_OUT8_Mp9@4989_g N_VDD_Mp9@4989_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4988 N_OUT9_Mp9@4988_d N_OUT8_Mp9@4988_g N_VDD_Mp9@4988_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4987 N_OUT9_Mn9@4987_d N_OUT8_Mn9@4987_g N_VSS_Mn9@4987_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4986 N_OUT9_Mn9@4986_d N_OUT8_Mn9@4986_g N_VSS_Mn9@4986_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4987 N_OUT9_Mp9@4987_d N_OUT8_Mp9@4987_g N_VDD_Mp9@4987_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4986 N_OUT9_Mp9@4986_d N_OUT8_Mp9@4986_g N_VDD_Mp9@4986_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4985 N_OUT9_Mn9@4985_d N_OUT8_Mn9@4985_g N_VSS_Mn9@4985_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4984 N_OUT9_Mn9@4984_d N_OUT8_Mn9@4984_g N_VSS_Mn9@4984_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4985 N_OUT9_Mp9@4985_d N_OUT8_Mp9@4985_g N_VDD_Mp9@4985_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4984 N_OUT9_Mp9@4984_d N_OUT8_Mp9@4984_g N_VDD_Mp9@4984_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4983 N_OUT9_Mn9@4983_d N_OUT8_Mn9@4983_g N_VSS_Mn9@4983_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4982 N_OUT9_Mn9@4982_d N_OUT8_Mn9@4982_g N_VSS_Mn9@4982_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4983 N_OUT9_Mp9@4983_d N_OUT8_Mp9@4983_g N_VDD_Mp9@4983_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4982 N_OUT9_Mp9@4982_d N_OUT8_Mp9@4982_g N_VDD_Mp9@4982_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4981 N_OUT9_Mn9@4981_d N_OUT8_Mn9@4981_g N_VSS_Mn9@4981_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4980 N_OUT9_Mn9@4980_d N_OUT8_Mn9@4980_g N_VSS_Mn9@4980_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4981 N_OUT9_Mp9@4981_d N_OUT8_Mp9@4981_g N_VDD_Mp9@4981_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4980 N_OUT9_Mp9@4980_d N_OUT8_Mp9@4980_g N_VDD_Mp9@4980_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4979 N_OUT9_Mn9@4979_d N_OUT8_Mn9@4979_g N_VSS_Mn9@4979_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4978 N_OUT9_Mn9@4978_d N_OUT8_Mn9@4978_g N_VSS_Mn9@4978_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4979 N_OUT9_Mp9@4979_d N_OUT8_Mp9@4979_g N_VDD_Mp9@4979_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4978 N_OUT9_Mp9@4978_d N_OUT8_Mp9@4978_g N_VDD_Mp9@4978_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4977 N_OUT9_Mn9@4977_d N_OUT8_Mn9@4977_g N_VSS_Mn9@4977_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4976 N_OUT9_Mn9@4976_d N_OUT8_Mn9@4976_g N_VSS_Mn9@4976_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4977 N_OUT9_Mp9@4977_d N_OUT8_Mp9@4977_g N_VDD_Mp9@4977_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4976 N_OUT9_Mp9@4976_d N_OUT8_Mp9@4976_g N_VDD_Mp9@4976_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4975 N_OUT9_Mn9@4975_d N_OUT8_Mn9@4975_g N_VSS_Mn9@4975_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4974 N_OUT9_Mn9@4974_d N_OUT8_Mn9@4974_g N_VSS_Mn9@4974_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4975 N_OUT9_Mp9@4975_d N_OUT8_Mp9@4975_g N_VDD_Mp9@4975_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4974 N_OUT9_Mp9@4974_d N_OUT8_Mp9@4974_g N_VDD_Mp9@4974_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4973 N_OUT9_Mn9@4973_d N_OUT8_Mn9@4973_g N_VSS_Mn9@4973_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4972 N_OUT9_Mn9@4972_d N_OUT8_Mn9@4972_g N_VSS_Mn9@4972_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4973 N_OUT9_Mp9@4973_d N_OUT8_Mp9@4973_g N_VDD_Mp9@4973_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4972 N_OUT9_Mp9@4972_d N_OUT8_Mp9@4972_g N_VDD_Mp9@4972_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4971 N_OUT9_Mn9@4971_d N_OUT8_Mn9@4971_g N_VSS_Mn9@4971_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4970 N_OUT9_Mn9@4970_d N_OUT8_Mn9@4970_g N_VSS_Mn9@4970_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4971 N_OUT9_Mp9@4971_d N_OUT8_Mp9@4971_g N_VDD_Mp9@4971_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4970 N_OUT9_Mp9@4970_d N_OUT8_Mp9@4970_g N_VDD_Mp9@4970_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4969 N_OUT9_Mn9@4969_d N_OUT8_Mn9@4969_g N_VSS_Mn9@4969_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4968 N_OUT9_Mn9@4968_d N_OUT8_Mn9@4968_g N_VSS_Mn9@4968_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4969 N_OUT9_Mp9@4969_d N_OUT8_Mp9@4969_g N_VDD_Mp9@4969_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4968 N_OUT9_Mp9@4968_d N_OUT8_Mp9@4968_g N_VDD_Mp9@4968_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4967 N_OUT9_Mn9@4967_d N_OUT8_Mn9@4967_g N_VSS_Mn9@4967_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4966 N_OUT9_Mn9@4966_d N_OUT8_Mn9@4966_g N_VSS_Mn9@4966_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4967 N_OUT9_Mp9@4967_d N_OUT8_Mp9@4967_g N_VDD_Mp9@4967_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4966 N_OUT9_Mp9@4966_d N_OUT8_Mp9@4966_g N_VDD_Mp9@4966_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4965 N_OUT9_Mn9@4965_d N_OUT8_Mn9@4965_g N_VSS_Mn9@4965_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4964 N_OUT9_Mn9@4964_d N_OUT8_Mn9@4964_g N_VSS_Mn9@4964_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4965 N_OUT9_Mp9@4965_d N_OUT8_Mp9@4965_g N_VDD_Mp9@4965_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4964 N_OUT9_Mp9@4964_d N_OUT8_Mp9@4964_g N_VDD_Mp9@4964_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4963 N_OUT9_Mn9@4963_d N_OUT8_Mn9@4963_g N_VSS_Mn9@4963_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4962 N_OUT9_Mn9@4962_d N_OUT8_Mn9@4962_g N_VSS_Mn9@4962_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4963 N_OUT9_Mp9@4963_d N_OUT8_Mp9@4963_g N_VDD_Mp9@4963_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4962 N_OUT9_Mp9@4962_d N_OUT8_Mp9@4962_g N_VDD_Mp9@4962_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4961 N_OUT9_Mn9@4961_d N_OUT8_Mn9@4961_g N_VSS_Mn9@4961_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4960 N_OUT9_Mn9@4960_d N_OUT8_Mn9@4960_g N_VSS_Mn9@4960_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4961 N_OUT9_Mp9@4961_d N_OUT8_Mp9@4961_g N_VDD_Mp9@4961_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4960 N_OUT9_Mp9@4960_d N_OUT8_Mp9@4960_g N_VDD_Mp9@4960_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4959 N_OUT9_Mn9@4959_d N_OUT8_Mn9@4959_g N_VSS_Mn9@4959_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4958 N_OUT9_Mn9@4958_d N_OUT8_Mn9@4958_g N_VSS_Mn9@4958_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4959 N_OUT9_Mp9@4959_d N_OUT8_Mp9@4959_g N_VDD_Mp9@4959_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4958 N_OUT9_Mp9@4958_d N_OUT8_Mp9@4958_g N_VDD_Mp9@4958_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4957 N_OUT9_Mn9@4957_d N_OUT8_Mn9@4957_g N_VSS_Mn9@4957_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4956 N_OUT9_Mn9@4956_d N_OUT8_Mn9@4956_g N_VSS_Mn9@4956_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4957 N_OUT9_Mp9@4957_d N_OUT8_Mp9@4957_g N_VDD_Mp9@4957_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4956 N_OUT9_Mp9@4956_d N_OUT8_Mp9@4956_g N_VDD_Mp9@4956_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4955 N_OUT9_Mn9@4955_d N_OUT8_Mn9@4955_g N_VSS_Mn9@4955_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4954 N_OUT9_Mn9@4954_d N_OUT8_Mn9@4954_g N_VSS_Mn9@4954_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4955 N_OUT9_Mp9@4955_d N_OUT8_Mp9@4955_g N_VDD_Mp9@4955_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4954 N_OUT9_Mp9@4954_d N_OUT8_Mp9@4954_g N_VDD_Mp9@4954_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4953 N_OUT9_Mn9@4953_d N_OUT8_Mn9@4953_g N_VSS_Mn9@4953_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4952 N_OUT9_Mn9@4952_d N_OUT8_Mn9@4952_g N_VSS_Mn9@4952_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4953 N_OUT9_Mp9@4953_d N_OUT8_Mp9@4953_g N_VDD_Mp9@4953_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4952 N_OUT9_Mp9@4952_d N_OUT8_Mp9@4952_g N_VDD_Mp9@4952_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4951 N_OUT9_Mn9@4951_d N_OUT8_Mn9@4951_g N_VSS_Mn9@4951_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4950 N_OUT9_Mn9@4950_d N_OUT8_Mn9@4950_g N_VSS_Mn9@4950_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4951 N_OUT9_Mp9@4951_d N_OUT8_Mp9@4951_g N_VDD_Mp9@4951_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4950 N_OUT9_Mp9@4950_d N_OUT8_Mp9@4950_g N_VDD_Mp9@4950_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4949 N_OUT9_Mn9@4949_d N_OUT8_Mn9@4949_g N_VSS_Mn9@4949_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4948 N_OUT9_Mn9@4948_d N_OUT8_Mn9@4948_g N_VSS_Mn9@4948_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4949 N_OUT9_Mp9@4949_d N_OUT8_Mp9@4949_g N_VDD_Mp9@4949_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4948 N_OUT9_Mp9@4948_d N_OUT8_Mp9@4948_g N_VDD_Mp9@4948_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4947 N_OUT9_Mn9@4947_d N_OUT8_Mn9@4947_g N_VSS_Mn9@4947_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4946 N_OUT9_Mn9@4946_d N_OUT8_Mn9@4946_g N_VSS_Mn9@4946_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4947 N_OUT9_Mp9@4947_d N_OUT8_Mp9@4947_g N_VDD_Mp9@4947_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4946 N_OUT9_Mp9@4946_d N_OUT8_Mp9@4946_g N_VDD_Mp9@4946_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4945 N_OUT9_Mn9@4945_d N_OUT8_Mn9@4945_g N_VSS_Mn9@4945_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4944 N_OUT9_Mn9@4944_d N_OUT8_Mn9@4944_g N_VSS_Mn9@4944_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4945 N_OUT9_Mp9@4945_d N_OUT8_Mp9@4945_g N_VDD_Mp9@4945_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4944 N_OUT9_Mp9@4944_d N_OUT8_Mp9@4944_g N_VDD_Mp9@4944_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4943 N_OUT9_Mn9@4943_d N_OUT8_Mn9@4943_g N_VSS_Mn9@4943_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4942 N_OUT9_Mn9@4942_d N_OUT8_Mn9@4942_g N_VSS_Mn9@4942_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4943 N_OUT9_Mp9@4943_d N_OUT8_Mp9@4943_g N_VDD_Mp9@4943_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4942 N_OUT9_Mp9@4942_d N_OUT8_Mp9@4942_g N_VDD_Mp9@4942_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4941 N_OUT9_Mn9@4941_d N_OUT8_Mn9@4941_g N_VSS_Mn9@4941_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4940 N_OUT9_Mn9@4940_d N_OUT8_Mn9@4940_g N_VSS_Mn9@4940_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4941 N_OUT9_Mp9@4941_d N_OUT8_Mp9@4941_g N_VDD_Mp9@4941_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4940 N_OUT9_Mp9@4940_d N_OUT8_Mp9@4940_g N_VDD_Mp9@4940_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4939 N_OUT9_Mn9@4939_d N_OUT8_Mn9@4939_g N_VSS_Mn9@4939_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4938 N_OUT9_Mn9@4938_d N_OUT8_Mn9@4938_g N_VSS_Mn9@4938_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4939 N_OUT9_Mp9@4939_d N_OUT8_Mp9@4939_g N_VDD_Mp9@4939_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4938 N_OUT9_Mp9@4938_d N_OUT8_Mp9@4938_g N_VDD_Mp9@4938_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4937 N_OUT9_Mn9@4937_d N_OUT8_Mn9@4937_g N_VSS_Mn9@4937_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4936 N_OUT9_Mn9@4936_d N_OUT8_Mn9@4936_g N_VSS_Mn9@4936_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4937 N_OUT9_Mp9@4937_d N_OUT8_Mp9@4937_g N_VDD_Mp9@4937_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4936 N_OUT9_Mp9@4936_d N_OUT8_Mp9@4936_g N_VDD_Mp9@4936_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4935 N_OUT9_Mn9@4935_d N_OUT8_Mn9@4935_g N_VSS_Mn9@4935_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4934 N_OUT9_Mn9@4934_d N_OUT8_Mn9@4934_g N_VSS_Mn9@4934_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4935 N_OUT9_Mp9@4935_d N_OUT8_Mp9@4935_g N_VDD_Mp9@4935_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4934 N_OUT9_Mp9@4934_d N_OUT8_Mp9@4934_g N_VDD_Mp9@4934_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4933 N_OUT9_Mn9@4933_d N_OUT8_Mn9@4933_g N_VSS_Mn9@4933_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4932 N_OUT9_Mn9@4932_d N_OUT8_Mn9@4932_g N_VSS_Mn9@4932_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4933 N_OUT9_Mp9@4933_d N_OUT8_Mp9@4933_g N_VDD_Mp9@4933_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4932 N_OUT9_Mp9@4932_d N_OUT8_Mp9@4932_g N_VDD_Mp9@4932_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4931 N_OUT9_Mn9@4931_d N_OUT8_Mn9@4931_g N_VSS_Mn9@4931_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4930 N_OUT9_Mn9@4930_d N_OUT8_Mn9@4930_g N_VSS_Mn9@4930_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4931 N_OUT9_Mp9@4931_d N_OUT8_Mp9@4931_g N_VDD_Mp9@4931_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4930 N_OUT9_Mp9@4930_d N_OUT8_Mp9@4930_g N_VDD_Mp9@4930_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4929 N_OUT9_Mn9@4929_d N_OUT8_Mn9@4929_g N_VSS_Mn9@4929_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4928 N_OUT9_Mn9@4928_d N_OUT8_Mn9@4928_g N_VSS_Mn9@4928_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4929 N_OUT9_Mp9@4929_d N_OUT8_Mp9@4929_g N_VDD_Mp9@4929_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4928 N_OUT9_Mp9@4928_d N_OUT8_Mp9@4928_g N_VDD_Mp9@4928_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4927 N_OUT9_Mn9@4927_d N_OUT8_Mn9@4927_g N_VSS_Mn9@4927_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4926 N_OUT9_Mn9@4926_d N_OUT8_Mn9@4926_g N_VSS_Mn9@4926_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4927 N_OUT9_Mp9@4927_d N_OUT8_Mp9@4927_g N_VDD_Mp9@4927_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4926 N_OUT9_Mp9@4926_d N_OUT8_Mp9@4926_g N_VDD_Mp9@4926_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4925 N_OUT9_Mn9@4925_d N_OUT8_Mn9@4925_g N_VSS_Mn9@4925_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4924 N_OUT9_Mn9@4924_d N_OUT8_Mn9@4924_g N_VSS_Mn9@4924_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4925 N_OUT9_Mp9@4925_d N_OUT8_Mp9@4925_g N_VDD_Mp9@4925_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4924 N_OUT9_Mp9@4924_d N_OUT8_Mp9@4924_g N_VDD_Mp9@4924_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4923 N_OUT9_Mn9@4923_d N_OUT8_Mn9@4923_g N_VSS_Mn9@4923_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4922 N_OUT9_Mn9@4922_d N_OUT8_Mn9@4922_g N_VSS_Mn9@4922_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4923 N_OUT9_Mp9@4923_d N_OUT8_Mp9@4923_g N_VDD_Mp9@4923_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4922 N_OUT9_Mp9@4922_d N_OUT8_Mp9@4922_g N_VDD_Mp9@4922_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4921 N_OUT9_Mn9@4921_d N_OUT8_Mn9@4921_g N_VSS_Mn9@4921_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4920 N_OUT9_Mn9@4920_d N_OUT8_Mn9@4920_g N_VSS_Mn9@4920_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4921 N_OUT9_Mp9@4921_d N_OUT8_Mp9@4921_g N_VDD_Mp9@4921_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4920 N_OUT9_Mp9@4920_d N_OUT8_Mp9@4920_g N_VDD_Mp9@4920_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4919 N_OUT9_Mn9@4919_d N_OUT8_Mn9@4919_g N_VSS_Mn9@4919_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4918 N_OUT9_Mn9@4918_d N_OUT8_Mn9@4918_g N_VSS_Mn9@4918_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4919 N_OUT9_Mp9@4919_d N_OUT8_Mp9@4919_g N_VDD_Mp9@4919_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4918 N_OUT9_Mp9@4918_d N_OUT8_Mp9@4918_g N_VDD_Mp9@4918_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4917 N_OUT9_Mn9@4917_d N_OUT8_Mn9@4917_g N_VSS_Mn9@4917_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4916 N_OUT9_Mn9@4916_d N_OUT8_Mn9@4916_g N_VSS_Mn9@4916_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4917 N_OUT9_Mp9@4917_d N_OUT8_Mp9@4917_g N_VDD_Mp9@4917_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4916 N_OUT9_Mp9@4916_d N_OUT8_Mp9@4916_g N_VDD_Mp9@4916_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4915 N_OUT9_Mn9@4915_d N_OUT8_Mn9@4915_g N_VSS_Mn9@4915_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4914 N_OUT9_Mn9@4914_d N_OUT8_Mn9@4914_g N_VSS_Mn9@4914_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4915 N_OUT9_Mp9@4915_d N_OUT8_Mp9@4915_g N_VDD_Mp9@4915_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4914 N_OUT9_Mp9@4914_d N_OUT8_Mp9@4914_g N_VDD_Mp9@4914_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4913 N_OUT9_Mn9@4913_d N_OUT8_Mn9@4913_g N_VSS_Mn9@4913_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4912 N_OUT9_Mn9@4912_d N_OUT8_Mn9@4912_g N_VSS_Mn9@4912_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4913 N_OUT9_Mp9@4913_d N_OUT8_Mp9@4913_g N_VDD_Mp9@4913_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4912 N_OUT9_Mp9@4912_d N_OUT8_Mp9@4912_g N_VDD_Mp9@4912_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4911 N_OUT9_Mn9@4911_d N_OUT8_Mn9@4911_g N_VSS_Mn9@4911_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4910 N_OUT9_Mn9@4910_d N_OUT8_Mn9@4910_g N_VSS_Mn9@4910_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4911 N_OUT9_Mp9@4911_d N_OUT8_Mp9@4911_g N_VDD_Mp9@4911_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4910 N_OUT9_Mp9@4910_d N_OUT8_Mp9@4910_g N_VDD_Mp9@4910_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4909 N_OUT9_Mn9@4909_d N_OUT8_Mn9@4909_g N_VSS_Mn9@4909_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4908 N_OUT9_Mn9@4908_d N_OUT8_Mn9@4908_g N_VSS_Mn9@4908_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4909 N_OUT9_Mp9@4909_d N_OUT8_Mp9@4909_g N_VDD_Mp9@4909_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4908 N_OUT9_Mp9@4908_d N_OUT8_Mp9@4908_g N_VDD_Mp9@4908_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4907 N_OUT9_Mn9@4907_d N_OUT8_Mn9@4907_g N_VSS_Mn9@4907_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4906 N_OUT9_Mn9@4906_d N_OUT8_Mn9@4906_g N_VSS_Mn9@4906_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4907 N_OUT9_Mp9@4907_d N_OUT8_Mp9@4907_g N_VDD_Mp9@4907_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4906 N_OUT9_Mp9@4906_d N_OUT8_Mp9@4906_g N_VDD_Mp9@4906_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4905 N_OUT9_Mn9@4905_d N_OUT8_Mn9@4905_g N_VSS_Mn9@4905_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4904 N_OUT9_Mn9@4904_d N_OUT8_Mn9@4904_g N_VSS_Mn9@4904_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4905 N_OUT9_Mp9@4905_d N_OUT8_Mp9@4905_g N_VDD_Mp9@4905_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4904 N_OUT9_Mp9@4904_d N_OUT8_Mp9@4904_g N_VDD_Mp9@4904_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4903 N_OUT9_Mn9@4903_d N_OUT8_Mn9@4903_g N_VSS_Mn9@4903_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4902 N_OUT9_Mn9@4902_d N_OUT8_Mn9@4902_g N_VSS_Mn9@4902_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4903 N_OUT9_Mp9@4903_d N_OUT8_Mp9@4903_g N_VDD_Mp9@4903_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4902 N_OUT9_Mp9@4902_d N_OUT8_Mp9@4902_g N_VDD_Mp9@4902_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4901 N_OUT9_Mn9@4901_d N_OUT8_Mn9@4901_g N_VSS_Mn9@4901_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4900 N_OUT9_Mn9@4900_d N_OUT8_Mn9@4900_g N_VSS_Mn9@4900_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4901 N_OUT9_Mp9@4901_d N_OUT8_Mp9@4901_g N_VDD_Mp9@4901_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4900 N_OUT9_Mp9@4900_d N_OUT8_Mp9@4900_g N_VDD_Mp9@4900_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4899 N_OUT9_Mn9@4899_d N_OUT8_Mn9@4899_g N_VSS_Mn9@4899_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4898 N_OUT9_Mn9@4898_d N_OUT8_Mn9@4898_g N_VSS_Mn9@4898_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4899 N_OUT9_Mp9@4899_d N_OUT8_Mp9@4899_g N_VDD_Mp9@4899_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4898 N_OUT9_Mp9@4898_d N_OUT8_Mp9@4898_g N_VDD_Mp9@4898_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4897 N_OUT9_Mn9@4897_d N_OUT8_Mn9@4897_g N_VSS_Mn9@4897_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4896 N_OUT9_Mn9@4896_d N_OUT8_Mn9@4896_g N_VSS_Mn9@4896_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4897 N_OUT9_Mp9@4897_d N_OUT8_Mp9@4897_g N_VDD_Mp9@4897_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4896 N_OUT9_Mp9@4896_d N_OUT8_Mp9@4896_g N_VDD_Mp9@4896_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4895 N_OUT9_Mn9@4895_d N_OUT8_Mn9@4895_g N_VSS_Mn9@4895_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4894 N_OUT9_Mn9@4894_d N_OUT8_Mn9@4894_g N_VSS_Mn9@4894_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4895 N_OUT9_Mp9@4895_d N_OUT8_Mp9@4895_g N_VDD_Mp9@4895_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4894 N_OUT9_Mp9@4894_d N_OUT8_Mp9@4894_g N_VDD_Mp9@4894_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4893 N_OUT9_Mn9@4893_d N_OUT8_Mn9@4893_g N_VSS_Mn9@4893_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4892 N_OUT9_Mn9@4892_d N_OUT8_Mn9@4892_g N_VSS_Mn9@4892_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4893 N_OUT9_Mp9@4893_d N_OUT8_Mp9@4893_g N_VDD_Mp9@4893_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4892 N_OUT9_Mp9@4892_d N_OUT8_Mp9@4892_g N_VDD_Mp9@4892_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4891 N_OUT9_Mn9@4891_d N_OUT8_Mn9@4891_g N_VSS_Mn9@4891_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4890 N_OUT9_Mn9@4890_d N_OUT8_Mn9@4890_g N_VSS_Mn9@4890_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4891 N_OUT9_Mp9@4891_d N_OUT8_Mp9@4891_g N_VDD_Mp9@4891_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4890 N_OUT9_Mp9@4890_d N_OUT8_Mp9@4890_g N_VDD_Mp9@4890_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4889 N_OUT9_Mn9@4889_d N_OUT8_Mn9@4889_g N_VSS_Mn9@4889_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4888 N_OUT9_Mn9@4888_d N_OUT8_Mn9@4888_g N_VSS_Mn9@4888_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4889 N_OUT9_Mp9@4889_d N_OUT8_Mp9@4889_g N_VDD_Mp9@4889_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4888 N_OUT9_Mp9@4888_d N_OUT8_Mp9@4888_g N_VDD_Mp9@4888_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4887 N_OUT9_Mn9@4887_d N_OUT8_Mn9@4887_g N_VSS_Mn9@4887_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4886 N_OUT9_Mn9@4886_d N_OUT8_Mn9@4886_g N_VSS_Mn9@4886_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4887 N_OUT9_Mp9@4887_d N_OUT8_Mp9@4887_g N_VDD_Mp9@4887_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4886 N_OUT9_Mp9@4886_d N_OUT8_Mp9@4886_g N_VDD_Mp9@4886_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4885 N_OUT9_Mn9@4885_d N_OUT8_Mn9@4885_g N_VSS_Mn9@4885_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4884 N_OUT9_Mn9@4884_d N_OUT8_Mn9@4884_g N_VSS_Mn9@4884_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4885 N_OUT9_Mp9@4885_d N_OUT8_Mp9@4885_g N_VDD_Mp9@4885_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4884 N_OUT9_Mp9@4884_d N_OUT8_Mp9@4884_g N_VDD_Mp9@4884_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4883 N_OUT9_Mn9@4883_d N_OUT8_Mn9@4883_g N_VSS_Mn9@4883_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4882 N_OUT9_Mn9@4882_d N_OUT8_Mn9@4882_g N_VSS_Mn9@4882_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4883 N_OUT9_Mp9@4883_d N_OUT8_Mp9@4883_g N_VDD_Mp9@4883_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4882 N_OUT9_Mp9@4882_d N_OUT8_Mp9@4882_g N_VDD_Mp9@4882_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4881 N_OUT9_Mn9@4881_d N_OUT8_Mn9@4881_g N_VSS_Mn9@4881_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4880 N_OUT9_Mn9@4880_d N_OUT8_Mn9@4880_g N_VSS_Mn9@4880_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4881 N_OUT9_Mp9@4881_d N_OUT8_Mp9@4881_g N_VDD_Mp9@4881_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4880 N_OUT9_Mp9@4880_d N_OUT8_Mp9@4880_g N_VDD_Mp9@4880_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4879 N_OUT9_Mn9@4879_d N_OUT8_Mn9@4879_g N_VSS_Mn9@4879_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4878 N_OUT9_Mn9@4878_d N_OUT8_Mn9@4878_g N_VSS_Mn9@4878_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4879 N_OUT9_Mp9@4879_d N_OUT8_Mp9@4879_g N_VDD_Mp9@4879_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4878 N_OUT9_Mp9@4878_d N_OUT8_Mp9@4878_g N_VDD_Mp9@4878_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4877 N_OUT9_Mn9@4877_d N_OUT8_Mn9@4877_g N_VSS_Mn9@4877_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4876 N_OUT9_Mn9@4876_d N_OUT8_Mn9@4876_g N_VSS_Mn9@4876_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4877 N_OUT9_Mp9@4877_d N_OUT8_Mp9@4877_g N_VDD_Mp9@4877_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4876 N_OUT9_Mp9@4876_d N_OUT8_Mp9@4876_g N_VDD_Mp9@4876_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4875 N_OUT9_Mn9@4875_d N_OUT8_Mn9@4875_g N_VSS_Mn9@4875_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4874 N_OUT9_Mn9@4874_d N_OUT8_Mn9@4874_g N_VSS_Mn9@4874_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4875 N_OUT9_Mp9@4875_d N_OUT8_Mp9@4875_g N_VDD_Mp9@4875_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4874 N_OUT9_Mp9@4874_d N_OUT8_Mp9@4874_g N_VDD_Mp9@4874_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4873 N_OUT9_Mn9@4873_d N_OUT8_Mn9@4873_g N_VSS_Mn9@4873_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4872 N_OUT9_Mn9@4872_d N_OUT8_Mn9@4872_g N_VSS_Mn9@4872_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4873 N_OUT9_Mp9@4873_d N_OUT8_Mp9@4873_g N_VDD_Mp9@4873_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4872 N_OUT9_Mp9@4872_d N_OUT8_Mp9@4872_g N_VDD_Mp9@4872_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4871 N_OUT9_Mn9@4871_d N_OUT8_Mn9@4871_g N_VSS_Mn9@4871_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4870 N_OUT9_Mn9@4870_d N_OUT8_Mn9@4870_g N_VSS_Mn9@4870_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4871 N_OUT9_Mp9@4871_d N_OUT8_Mp9@4871_g N_VDD_Mp9@4871_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4870 N_OUT9_Mp9@4870_d N_OUT8_Mp9@4870_g N_VDD_Mp9@4870_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4869 N_OUT9_Mn9@4869_d N_OUT8_Mn9@4869_g N_VSS_Mn9@4869_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4868 N_OUT9_Mn9@4868_d N_OUT8_Mn9@4868_g N_VSS_Mn9@4868_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4869 N_OUT9_Mp9@4869_d N_OUT8_Mp9@4869_g N_VDD_Mp9@4869_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4868 N_OUT9_Mp9@4868_d N_OUT8_Mp9@4868_g N_VDD_Mp9@4868_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4867 N_OUT9_Mn9@4867_d N_OUT8_Mn9@4867_g N_VSS_Mn9@4867_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4866 N_OUT9_Mn9@4866_d N_OUT8_Mn9@4866_g N_VSS_Mn9@4866_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4867 N_OUT9_Mp9@4867_d N_OUT8_Mp9@4867_g N_VDD_Mp9@4867_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4866 N_OUT9_Mp9@4866_d N_OUT8_Mp9@4866_g N_VDD_Mp9@4866_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4865 N_OUT9_Mn9@4865_d N_OUT8_Mn9@4865_g N_VSS_Mn9@4865_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4864 N_OUT9_Mn9@4864_d N_OUT8_Mn9@4864_g N_VSS_Mn9@4864_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4865 N_OUT9_Mp9@4865_d N_OUT8_Mp9@4865_g N_VDD_Mp9@4865_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4864 N_OUT9_Mp9@4864_d N_OUT8_Mp9@4864_g N_VDD_Mp9@4864_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4863 N_OUT9_Mn9@4863_d N_OUT8_Mn9@4863_g N_VSS_Mn9@4863_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4862 N_OUT9_Mn9@4862_d N_OUT8_Mn9@4862_g N_VSS_Mn9@4862_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4863 N_OUT9_Mp9@4863_d N_OUT8_Mp9@4863_g N_VDD_Mp9@4863_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4862 N_OUT9_Mp9@4862_d N_OUT8_Mp9@4862_g N_VDD_Mp9@4862_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4861 N_OUT9_Mn9@4861_d N_OUT8_Mn9@4861_g N_VSS_Mn9@4861_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4860 N_OUT9_Mn9@4860_d N_OUT8_Mn9@4860_g N_VSS_Mn9@4860_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4861 N_OUT9_Mp9@4861_d N_OUT8_Mp9@4861_g N_VDD_Mp9@4861_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4860 N_OUT9_Mp9@4860_d N_OUT8_Mp9@4860_g N_VDD_Mp9@4860_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4859 N_OUT9_Mn9@4859_d N_OUT8_Mn9@4859_g N_VSS_Mn9@4859_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4858 N_OUT9_Mn9@4858_d N_OUT8_Mn9@4858_g N_VSS_Mn9@4858_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4859 N_OUT9_Mp9@4859_d N_OUT8_Mp9@4859_g N_VDD_Mp9@4859_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4858 N_OUT9_Mp9@4858_d N_OUT8_Mp9@4858_g N_VDD_Mp9@4858_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4857 N_OUT9_Mn9@4857_d N_OUT8_Mn9@4857_g N_VSS_Mn9@4857_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4856 N_OUT9_Mn9@4856_d N_OUT8_Mn9@4856_g N_VSS_Mn9@4856_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4857 N_OUT9_Mp9@4857_d N_OUT8_Mp9@4857_g N_VDD_Mp9@4857_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4856 N_OUT9_Mp9@4856_d N_OUT8_Mp9@4856_g N_VDD_Mp9@4856_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4855 N_OUT9_Mn9@4855_d N_OUT8_Mn9@4855_g N_VSS_Mn9@4855_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4854 N_OUT9_Mn9@4854_d N_OUT8_Mn9@4854_g N_VSS_Mn9@4854_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4855 N_OUT9_Mp9@4855_d N_OUT8_Mp9@4855_g N_VDD_Mp9@4855_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4854 N_OUT9_Mp9@4854_d N_OUT8_Mp9@4854_g N_VDD_Mp9@4854_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4853 N_OUT9_Mn9@4853_d N_OUT8_Mn9@4853_g N_VSS_Mn9@4853_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4852 N_OUT9_Mn9@4852_d N_OUT8_Mn9@4852_g N_VSS_Mn9@4852_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4853 N_OUT9_Mp9@4853_d N_OUT8_Mp9@4853_g N_VDD_Mp9@4853_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4852 N_OUT9_Mp9@4852_d N_OUT8_Mp9@4852_g N_VDD_Mp9@4852_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4851 N_OUT9_Mn9@4851_d N_OUT8_Mn9@4851_g N_VSS_Mn9@4851_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4850 N_OUT9_Mn9@4850_d N_OUT8_Mn9@4850_g N_VSS_Mn9@4850_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4851 N_OUT9_Mp9@4851_d N_OUT8_Mp9@4851_g N_VDD_Mp9@4851_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4850 N_OUT9_Mp9@4850_d N_OUT8_Mp9@4850_g N_VDD_Mp9@4850_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4849 N_OUT9_Mn9@4849_d N_OUT8_Mn9@4849_g N_VSS_Mn9@4849_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4848 N_OUT9_Mn9@4848_d N_OUT8_Mn9@4848_g N_VSS_Mn9@4848_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4849 N_OUT9_Mp9@4849_d N_OUT8_Mp9@4849_g N_VDD_Mp9@4849_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4848 N_OUT9_Mp9@4848_d N_OUT8_Mp9@4848_g N_VDD_Mp9@4848_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4847 N_OUT9_Mn9@4847_d N_OUT8_Mn9@4847_g N_VSS_Mn9@4847_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4846 N_OUT9_Mn9@4846_d N_OUT8_Mn9@4846_g N_VSS_Mn9@4846_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4847 N_OUT9_Mp9@4847_d N_OUT8_Mp9@4847_g N_VDD_Mp9@4847_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4846 N_OUT9_Mp9@4846_d N_OUT8_Mp9@4846_g N_VDD_Mp9@4846_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4845 N_OUT9_Mn9@4845_d N_OUT8_Mn9@4845_g N_VSS_Mn9@4845_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4844 N_OUT9_Mn9@4844_d N_OUT8_Mn9@4844_g N_VSS_Mn9@4844_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4845 N_OUT9_Mp9@4845_d N_OUT8_Mp9@4845_g N_VDD_Mp9@4845_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4844 N_OUT9_Mp9@4844_d N_OUT8_Mp9@4844_g N_VDD_Mp9@4844_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4843 N_OUT9_Mn9@4843_d N_OUT8_Mn9@4843_g N_VSS_Mn9@4843_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4842 N_OUT9_Mn9@4842_d N_OUT8_Mn9@4842_g N_VSS_Mn9@4842_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4843 N_OUT9_Mp9@4843_d N_OUT8_Mp9@4843_g N_VDD_Mp9@4843_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4842 N_OUT9_Mp9@4842_d N_OUT8_Mp9@4842_g N_VDD_Mp9@4842_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4841 N_OUT9_Mn9@4841_d N_OUT8_Mn9@4841_g N_VSS_Mn9@4841_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4840 N_OUT9_Mn9@4840_d N_OUT8_Mn9@4840_g N_VSS_Mn9@4840_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4841 N_OUT9_Mp9@4841_d N_OUT8_Mp9@4841_g N_VDD_Mp9@4841_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4840 N_OUT9_Mp9@4840_d N_OUT8_Mp9@4840_g N_VDD_Mp9@4840_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4839 N_OUT9_Mn9@4839_d N_OUT8_Mn9@4839_g N_VSS_Mn9@4839_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4838 N_OUT9_Mn9@4838_d N_OUT8_Mn9@4838_g N_VSS_Mn9@4838_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4839 N_OUT9_Mp9@4839_d N_OUT8_Mp9@4839_g N_VDD_Mp9@4839_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4838 N_OUT9_Mp9@4838_d N_OUT8_Mp9@4838_g N_VDD_Mp9@4838_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4837 N_OUT9_Mn9@4837_d N_OUT8_Mn9@4837_g N_VSS_Mn9@4837_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4836 N_OUT9_Mn9@4836_d N_OUT8_Mn9@4836_g N_VSS_Mn9@4836_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4837 N_OUT9_Mp9@4837_d N_OUT8_Mp9@4837_g N_VDD_Mp9@4837_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4836 N_OUT9_Mp9@4836_d N_OUT8_Mp9@4836_g N_VDD_Mp9@4836_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4835 N_OUT9_Mn9@4835_d N_OUT8_Mn9@4835_g N_VSS_Mn9@4835_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4834 N_OUT9_Mn9@4834_d N_OUT8_Mn9@4834_g N_VSS_Mn9@4834_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4835 N_OUT9_Mp9@4835_d N_OUT8_Mp9@4835_g N_VDD_Mp9@4835_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4834 N_OUT9_Mp9@4834_d N_OUT8_Mp9@4834_g N_VDD_Mp9@4834_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4833 N_OUT9_Mn9@4833_d N_OUT8_Mn9@4833_g N_VSS_Mn9@4833_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4832 N_OUT9_Mn9@4832_d N_OUT8_Mn9@4832_g N_VSS_Mn9@4832_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4833 N_OUT9_Mp9@4833_d N_OUT8_Mp9@4833_g N_VDD_Mp9@4833_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4832 N_OUT9_Mp9@4832_d N_OUT8_Mp9@4832_g N_VDD_Mp9@4832_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4831 N_OUT9_Mn9@4831_d N_OUT8_Mn9@4831_g N_VSS_Mn9@4831_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4830 N_OUT9_Mn9@4830_d N_OUT8_Mn9@4830_g N_VSS_Mn9@4830_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4831 N_OUT9_Mp9@4831_d N_OUT8_Mp9@4831_g N_VDD_Mp9@4831_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4830 N_OUT9_Mp9@4830_d N_OUT8_Mp9@4830_g N_VDD_Mp9@4830_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4829 N_OUT9_Mn9@4829_d N_OUT8_Mn9@4829_g N_VSS_Mn9@4829_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4828 N_OUT9_Mn9@4828_d N_OUT8_Mn9@4828_g N_VSS_Mn9@4828_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4829 N_OUT9_Mp9@4829_d N_OUT8_Mp9@4829_g N_VDD_Mp9@4829_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4828 N_OUT9_Mp9@4828_d N_OUT8_Mp9@4828_g N_VDD_Mp9@4828_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4827 N_OUT9_Mn9@4827_d N_OUT8_Mn9@4827_g N_VSS_Mn9@4827_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4826 N_OUT9_Mn9@4826_d N_OUT8_Mn9@4826_g N_VSS_Mn9@4826_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4827 N_OUT9_Mp9@4827_d N_OUT8_Mp9@4827_g N_VDD_Mp9@4827_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4826 N_OUT9_Mp9@4826_d N_OUT8_Mp9@4826_g N_VDD_Mp9@4826_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4825 N_OUT9_Mn9@4825_d N_OUT8_Mn9@4825_g N_VSS_Mn9@4825_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4824 N_OUT9_Mn9@4824_d N_OUT8_Mn9@4824_g N_VSS_Mn9@4824_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4825 N_OUT9_Mp9@4825_d N_OUT8_Mp9@4825_g N_VDD_Mp9@4825_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4824 N_OUT9_Mp9@4824_d N_OUT8_Mp9@4824_g N_VDD_Mp9@4824_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4823 N_OUT9_Mn9@4823_d N_OUT8_Mn9@4823_g N_VSS_Mn9@4823_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4822 N_OUT9_Mn9@4822_d N_OUT8_Mn9@4822_g N_VSS_Mn9@4822_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4823 N_OUT9_Mp9@4823_d N_OUT8_Mp9@4823_g N_VDD_Mp9@4823_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4822 N_OUT9_Mp9@4822_d N_OUT8_Mp9@4822_g N_VDD_Mp9@4822_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4821 N_OUT9_Mn9@4821_d N_OUT8_Mn9@4821_g N_VSS_Mn9@4821_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4820 N_OUT9_Mn9@4820_d N_OUT8_Mn9@4820_g N_VSS_Mn9@4820_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4821 N_OUT9_Mp9@4821_d N_OUT8_Mp9@4821_g N_VDD_Mp9@4821_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4820 N_OUT9_Mp9@4820_d N_OUT8_Mp9@4820_g N_VDD_Mp9@4820_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4819 N_OUT9_Mn9@4819_d N_OUT8_Mn9@4819_g N_VSS_Mn9@4819_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4818 N_OUT9_Mn9@4818_d N_OUT8_Mn9@4818_g N_VSS_Mn9@4818_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4819 N_OUT9_Mp9@4819_d N_OUT8_Mp9@4819_g N_VDD_Mp9@4819_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4818 N_OUT9_Mp9@4818_d N_OUT8_Mp9@4818_g N_VDD_Mp9@4818_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4817 N_OUT9_Mn9@4817_d N_OUT8_Mn9@4817_g N_VSS_Mn9@4817_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4816 N_OUT9_Mn9@4816_d N_OUT8_Mn9@4816_g N_VSS_Mn9@4816_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4817 N_OUT9_Mp9@4817_d N_OUT8_Mp9@4817_g N_VDD_Mp9@4817_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4816 N_OUT9_Mp9@4816_d N_OUT8_Mp9@4816_g N_VDD_Mp9@4816_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4815 N_OUT9_Mn9@4815_d N_OUT8_Mn9@4815_g N_VSS_Mn9@4815_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4814 N_OUT9_Mn9@4814_d N_OUT8_Mn9@4814_g N_VSS_Mn9@4814_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4815 N_OUT9_Mp9@4815_d N_OUT8_Mp9@4815_g N_VDD_Mp9@4815_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4814 N_OUT9_Mp9@4814_d N_OUT8_Mp9@4814_g N_VDD_Mp9@4814_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4813 N_OUT9_Mn9@4813_d N_OUT8_Mn9@4813_g N_VSS_Mn9@4813_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4812 N_OUT9_Mn9@4812_d N_OUT8_Mn9@4812_g N_VSS_Mn9@4812_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4813 N_OUT9_Mp9@4813_d N_OUT8_Mp9@4813_g N_VDD_Mp9@4813_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4812 N_OUT9_Mp9@4812_d N_OUT8_Mp9@4812_g N_VDD_Mp9@4812_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4811 N_OUT9_Mn9@4811_d N_OUT8_Mn9@4811_g N_VSS_Mn9@4811_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4810 N_OUT9_Mn9@4810_d N_OUT8_Mn9@4810_g N_VSS_Mn9@4810_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4811 N_OUT9_Mp9@4811_d N_OUT8_Mp9@4811_g N_VDD_Mp9@4811_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4810 N_OUT9_Mp9@4810_d N_OUT8_Mp9@4810_g N_VDD_Mp9@4810_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4809 N_OUT9_Mn9@4809_d N_OUT8_Mn9@4809_g N_VSS_Mn9@4809_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4808 N_OUT9_Mn9@4808_d N_OUT8_Mn9@4808_g N_VSS_Mn9@4808_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4809 N_OUT9_Mp9@4809_d N_OUT8_Mp9@4809_g N_VDD_Mp9@4809_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4808 N_OUT9_Mp9@4808_d N_OUT8_Mp9@4808_g N_VDD_Mp9@4808_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4807 N_OUT9_Mn9@4807_d N_OUT8_Mn9@4807_g N_VSS_Mn9@4807_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4806 N_OUT9_Mn9@4806_d N_OUT8_Mn9@4806_g N_VSS_Mn9@4806_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4807 N_OUT9_Mp9@4807_d N_OUT8_Mp9@4807_g N_VDD_Mp9@4807_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4806 N_OUT9_Mp9@4806_d N_OUT8_Mp9@4806_g N_VDD_Mp9@4806_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4805 N_OUT9_Mn9@4805_d N_OUT8_Mn9@4805_g N_VSS_Mn9@4805_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4804 N_OUT9_Mn9@4804_d N_OUT8_Mn9@4804_g N_VSS_Mn9@4804_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4805 N_OUT9_Mp9@4805_d N_OUT8_Mp9@4805_g N_VDD_Mp9@4805_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4804 N_OUT9_Mp9@4804_d N_OUT8_Mp9@4804_g N_VDD_Mp9@4804_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4803 N_OUT9_Mn9@4803_d N_OUT8_Mn9@4803_g N_VSS_Mn9@4803_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4802 N_OUT9_Mn9@4802_d N_OUT8_Mn9@4802_g N_VSS_Mn9@4802_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4803 N_OUT9_Mp9@4803_d N_OUT8_Mp9@4803_g N_VDD_Mp9@4803_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4802 N_OUT9_Mp9@4802_d N_OUT8_Mp9@4802_g N_VDD_Mp9@4802_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4801 N_OUT9_Mn9@4801_d N_OUT8_Mn9@4801_g N_VSS_Mn9@4801_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4800 N_OUT9_Mn9@4800_d N_OUT8_Mn9@4800_g N_VSS_Mn9@4800_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4801 N_OUT9_Mp9@4801_d N_OUT8_Mp9@4801_g N_VDD_Mp9@4801_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4800 N_OUT9_Mp9@4800_d N_OUT8_Mp9@4800_g N_VDD_Mp9@4800_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4799 N_OUT9_Mn9@4799_d N_OUT8_Mn9@4799_g N_VSS_Mn9@4799_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4798 N_OUT9_Mn9@4798_d N_OUT8_Mn9@4798_g N_VSS_Mn9@4798_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4799 N_OUT9_Mp9@4799_d N_OUT8_Mp9@4799_g N_VDD_Mp9@4799_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4798 N_OUT9_Mp9@4798_d N_OUT8_Mp9@4798_g N_VDD_Mp9@4798_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4797 N_OUT9_Mn9@4797_d N_OUT8_Mn9@4797_g N_VSS_Mn9@4797_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4796 N_OUT9_Mn9@4796_d N_OUT8_Mn9@4796_g N_VSS_Mn9@4796_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4797 N_OUT9_Mp9@4797_d N_OUT8_Mp9@4797_g N_VDD_Mp9@4797_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4796 N_OUT9_Mp9@4796_d N_OUT8_Mp9@4796_g N_VDD_Mp9@4796_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4795 N_OUT9_Mn9@4795_d N_OUT8_Mn9@4795_g N_VSS_Mn9@4795_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4794 N_OUT9_Mn9@4794_d N_OUT8_Mn9@4794_g N_VSS_Mn9@4794_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4795 N_OUT9_Mp9@4795_d N_OUT8_Mp9@4795_g N_VDD_Mp9@4795_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4794 N_OUT9_Mp9@4794_d N_OUT8_Mp9@4794_g N_VDD_Mp9@4794_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4793 N_OUT9_Mn9@4793_d N_OUT8_Mn9@4793_g N_VSS_Mn9@4793_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4792 N_OUT9_Mn9@4792_d N_OUT8_Mn9@4792_g N_VSS_Mn9@4792_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4793 N_OUT9_Mp9@4793_d N_OUT8_Mp9@4793_g N_VDD_Mp9@4793_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4792 N_OUT9_Mp9@4792_d N_OUT8_Mp9@4792_g N_VDD_Mp9@4792_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4791 N_OUT9_Mn9@4791_d N_OUT8_Mn9@4791_g N_VSS_Mn9@4791_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4790 N_OUT9_Mn9@4790_d N_OUT8_Mn9@4790_g N_VSS_Mn9@4790_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4791 N_OUT9_Mp9@4791_d N_OUT8_Mp9@4791_g N_VDD_Mp9@4791_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4790 N_OUT9_Mp9@4790_d N_OUT8_Mp9@4790_g N_VDD_Mp9@4790_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4789 N_OUT9_Mn9@4789_d N_OUT8_Mn9@4789_g N_VSS_Mn9@4789_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4788 N_OUT9_Mn9@4788_d N_OUT8_Mn9@4788_g N_VSS_Mn9@4788_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4789 N_OUT9_Mp9@4789_d N_OUT8_Mp9@4789_g N_VDD_Mp9@4789_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4788 N_OUT9_Mp9@4788_d N_OUT8_Mp9@4788_g N_VDD_Mp9@4788_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4787 N_OUT9_Mn9@4787_d N_OUT8_Mn9@4787_g N_VSS_Mn9@4787_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4786 N_OUT9_Mn9@4786_d N_OUT8_Mn9@4786_g N_VSS_Mn9@4786_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4787 N_OUT9_Mp9@4787_d N_OUT8_Mp9@4787_g N_VDD_Mp9@4787_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4786 N_OUT9_Mp9@4786_d N_OUT8_Mp9@4786_g N_VDD_Mp9@4786_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4785 N_OUT9_Mn9@4785_d N_OUT8_Mn9@4785_g N_VSS_Mn9@4785_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4784 N_OUT9_Mn9@4784_d N_OUT8_Mn9@4784_g N_VSS_Mn9@4784_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4785 N_OUT9_Mp9@4785_d N_OUT8_Mp9@4785_g N_VDD_Mp9@4785_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4784 N_OUT9_Mp9@4784_d N_OUT8_Mp9@4784_g N_VDD_Mp9@4784_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4783 N_OUT9_Mn9@4783_d N_OUT8_Mn9@4783_g N_VSS_Mn9@4783_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4782 N_OUT9_Mn9@4782_d N_OUT8_Mn9@4782_g N_VSS_Mn9@4782_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4783 N_OUT9_Mp9@4783_d N_OUT8_Mp9@4783_g N_VDD_Mp9@4783_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4782 N_OUT9_Mp9@4782_d N_OUT8_Mp9@4782_g N_VDD_Mp9@4782_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4781 N_OUT9_Mn9@4781_d N_OUT8_Mn9@4781_g N_VSS_Mn9@4781_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4780 N_OUT9_Mn9@4780_d N_OUT8_Mn9@4780_g N_VSS_Mn9@4780_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4781 N_OUT9_Mp9@4781_d N_OUT8_Mp9@4781_g N_VDD_Mp9@4781_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4780 N_OUT9_Mp9@4780_d N_OUT8_Mp9@4780_g N_VDD_Mp9@4780_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4779 N_OUT9_Mn9@4779_d N_OUT8_Mn9@4779_g N_VSS_Mn9@4779_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4778 N_OUT9_Mn9@4778_d N_OUT8_Mn9@4778_g N_VSS_Mn9@4778_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4779 N_OUT9_Mp9@4779_d N_OUT8_Mp9@4779_g N_VDD_Mp9@4779_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4778 N_OUT9_Mp9@4778_d N_OUT8_Mp9@4778_g N_VDD_Mp9@4778_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4777 N_OUT9_Mn9@4777_d N_OUT8_Mn9@4777_g N_VSS_Mn9@4777_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4776 N_OUT9_Mn9@4776_d N_OUT8_Mn9@4776_g N_VSS_Mn9@4776_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4777 N_OUT9_Mp9@4777_d N_OUT8_Mp9@4777_g N_VDD_Mp9@4777_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4776 N_OUT9_Mp9@4776_d N_OUT8_Mp9@4776_g N_VDD_Mp9@4776_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4775 N_OUT9_Mn9@4775_d N_OUT8_Mn9@4775_g N_VSS_Mn9@4775_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4774 N_OUT9_Mn9@4774_d N_OUT8_Mn9@4774_g N_VSS_Mn9@4774_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4775 N_OUT9_Mp9@4775_d N_OUT8_Mp9@4775_g N_VDD_Mp9@4775_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4774 N_OUT9_Mp9@4774_d N_OUT8_Mp9@4774_g N_VDD_Mp9@4774_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4773 N_OUT9_Mn9@4773_d N_OUT8_Mn9@4773_g N_VSS_Mn9@4773_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4772 N_OUT9_Mn9@4772_d N_OUT8_Mn9@4772_g N_VSS_Mn9@4772_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4773 N_OUT9_Mp9@4773_d N_OUT8_Mp9@4773_g N_VDD_Mp9@4773_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4772 N_OUT9_Mp9@4772_d N_OUT8_Mp9@4772_g N_VDD_Mp9@4772_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4771 N_OUT9_Mn9@4771_d N_OUT8_Mn9@4771_g N_VSS_Mn9@4771_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4770 N_OUT9_Mn9@4770_d N_OUT8_Mn9@4770_g N_VSS_Mn9@4770_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4771 N_OUT9_Mp9@4771_d N_OUT8_Mp9@4771_g N_VDD_Mp9@4771_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4770 N_OUT9_Mp9@4770_d N_OUT8_Mp9@4770_g N_VDD_Mp9@4770_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4769 N_OUT9_Mn9@4769_d N_OUT8_Mn9@4769_g N_VSS_Mn9@4769_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4768 N_OUT9_Mn9@4768_d N_OUT8_Mn9@4768_g N_VSS_Mn9@4768_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4769 N_OUT9_Mp9@4769_d N_OUT8_Mp9@4769_g N_VDD_Mp9@4769_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4768 N_OUT9_Mp9@4768_d N_OUT8_Mp9@4768_g N_VDD_Mp9@4768_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4767 N_OUT9_Mn9@4767_d N_OUT8_Mn9@4767_g N_VSS_Mn9@4767_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4766 N_OUT9_Mn9@4766_d N_OUT8_Mn9@4766_g N_VSS_Mn9@4766_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4767 N_OUT9_Mp9@4767_d N_OUT8_Mp9@4767_g N_VDD_Mp9@4767_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4766 N_OUT9_Mp9@4766_d N_OUT8_Mp9@4766_g N_VDD_Mp9@4766_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4765 N_OUT9_Mn9@4765_d N_OUT8_Mn9@4765_g N_VSS_Mn9@4765_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4764 N_OUT9_Mn9@4764_d N_OUT8_Mn9@4764_g N_VSS_Mn9@4764_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4765 N_OUT9_Mp9@4765_d N_OUT8_Mp9@4765_g N_VDD_Mp9@4765_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4764 N_OUT9_Mp9@4764_d N_OUT8_Mp9@4764_g N_VDD_Mp9@4764_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4763 N_OUT9_Mn9@4763_d N_OUT8_Mn9@4763_g N_VSS_Mn9@4763_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4762 N_OUT9_Mn9@4762_d N_OUT8_Mn9@4762_g N_VSS_Mn9@4762_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4763 N_OUT9_Mp9@4763_d N_OUT8_Mp9@4763_g N_VDD_Mp9@4763_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4762 N_OUT9_Mp9@4762_d N_OUT8_Mp9@4762_g N_VDD_Mp9@4762_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4761 N_OUT9_Mn9@4761_d N_OUT8_Mn9@4761_g N_VSS_Mn9@4761_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4760 N_OUT9_Mn9@4760_d N_OUT8_Mn9@4760_g N_VSS_Mn9@4760_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4761 N_OUT9_Mp9@4761_d N_OUT8_Mp9@4761_g N_VDD_Mp9@4761_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4760 N_OUT9_Mp9@4760_d N_OUT8_Mp9@4760_g N_VDD_Mp9@4760_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4759 N_OUT9_Mn9@4759_d N_OUT8_Mn9@4759_g N_VSS_Mn9@4759_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4758 N_OUT9_Mn9@4758_d N_OUT8_Mn9@4758_g N_VSS_Mn9@4758_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4759 N_OUT9_Mp9@4759_d N_OUT8_Mp9@4759_g N_VDD_Mp9@4759_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4758 N_OUT9_Mp9@4758_d N_OUT8_Mp9@4758_g N_VDD_Mp9@4758_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4757 N_OUT9_Mn9@4757_d N_OUT8_Mn9@4757_g N_VSS_Mn9@4757_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4756 N_OUT9_Mn9@4756_d N_OUT8_Mn9@4756_g N_VSS_Mn9@4756_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4757 N_OUT9_Mp9@4757_d N_OUT8_Mp9@4757_g N_VDD_Mp9@4757_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4756 N_OUT9_Mp9@4756_d N_OUT8_Mp9@4756_g N_VDD_Mp9@4756_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4755 N_OUT9_Mn9@4755_d N_OUT8_Mn9@4755_g N_VSS_Mn9@4755_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4754 N_OUT9_Mn9@4754_d N_OUT8_Mn9@4754_g N_VSS_Mn9@4754_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4755 N_OUT9_Mp9@4755_d N_OUT8_Mp9@4755_g N_VDD_Mp9@4755_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4754 N_OUT9_Mp9@4754_d N_OUT8_Mp9@4754_g N_VDD_Mp9@4754_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4753 N_OUT9_Mn9@4753_d N_OUT8_Mn9@4753_g N_VSS_Mn9@4753_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4752 N_OUT9_Mn9@4752_d N_OUT8_Mn9@4752_g N_VSS_Mn9@4752_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4753 N_OUT9_Mp9@4753_d N_OUT8_Mp9@4753_g N_VDD_Mp9@4753_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4752 N_OUT9_Mp9@4752_d N_OUT8_Mp9@4752_g N_VDD_Mp9@4752_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4751 N_OUT9_Mn9@4751_d N_OUT8_Mn9@4751_g N_VSS_Mn9@4751_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4750 N_OUT9_Mn9@4750_d N_OUT8_Mn9@4750_g N_VSS_Mn9@4750_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4751 N_OUT9_Mp9@4751_d N_OUT8_Mp9@4751_g N_VDD_Mp9@4751_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4750 N_OUT9_Mp9@4750_d N_OUT8_Mp9@4750_g N_VDD_Mp9@4750_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4749 N_OUT9_Mn9@4749_d N_OUT8_Mn9@4749_g N_VSS_Mn9@4749_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4748 N_OUT9_Mn9@4748_d N_OUT8_Mn9@4748_g N_VSS_Mn9@4748_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4749 N_OUT9_Mp9@4749_d N_OUT8_Mp9@4749_g N_VDD_Mp9@4749_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4748 N_OUT9_Mp9@4748_d N_OUT8_Mp9@4748_g N_VDD_Mp9@4748_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4747 N_OUT9_Mn9@4747_d N_OUT8_Mn9@4747_g N_VSS_Mn9@4747_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4746 N_OUT9_Mn9@4746_d N_OUT8_Mn9@4746_g N_VSS_Mn9@4746_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4747 N_OUT9_Mp9@4747_d N_OUT8_Mp9@4747_g N_VDD_Mp9@4747_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4746 N_OUT9_Mp9@4746_d N_OUT8_Mp9@4746_g N_VDD_Mp9@4746_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4745 N_OUT9_Mn9@4745_d N_OUT8_Mn9@4745_g N_VSS_Mn9@4745_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4744 N_OUT9_Mn9@4744_d N_OUT8_Mn9@4744_g N_VSS_Mn9@4744_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4745 N_OUT9_Mp9@4745_d N_OUT8_Mp9@4745_g N_VDD_Mp9@4745_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4744 N_OUT9_Mp9@4744_d N_OUT8_Mp9@4744_g N_VDD_Mp9@4744_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4743 N_OUT9_Mn9@4743_d N_OUT8_Mn9@4743_g N_VSS_Mn9@4743_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4742 N_OUT9_Mn9@4742_d N_OUT8_Mn9@4742_g N_VSS_Mn9@4742_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4743 N_OUT9_Mp9@4743_d N_OUT8_Mp9@4743_g N_VDD_Mp9@4743_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4742 N_OUT9_Mp9@4742_d N_OUT8_Mp9@4742_g N_VDD_Mp9@4742_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4741 N_OUT9_Mn9@4741_d N_OUT8_Mn9@4741_g N_VSS_Mn9@4741_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4740 N_OUT9_Mn9@4740_d N_OUT8_Mn9@4740_g N_VSS_Mn9@4740_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4741 N_OUT9_Mp9@4741_d N_OUT8_Mp9@4741_g N_VDD_Mp9@4741_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4740 N_OUT9_Mp9@4740_d N_OUT8_Mp9@4740_g N_VDD_Mp9@4740_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4739 N_OUT9_Mn9@4739_d N_OUT8_Mn9@4739_g N_VSS_Mn9@4739_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4738 N_OUT9_Mn9@4738_d N_OUT8_Mn9@4738_g N_VSS_Mn9@4738_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4739 N_OUT9_Mp9@4739_d N_OUT8_Mp9@4739_g N_VDD_Mp9@4739_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4738 N_OUT9_Mp9@4738_d N_OUT8_Mp9@4738_g N_VDD_Mp9@4738_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4737 N_OUT9_Mn9@4737_d N_OUT8_Mn9@4737_g N_VSS_Mn9@4737_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4736 N_OUT9_Mn9@4736_d N_OUT8_Mn9@4736_g N_VSS_Mn9@4736_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4737 N_OUT9_Mp9@4737_d N_OUT8_Mp9@4737_g N_VDD_Mp9@4737_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4736 N_OUT9_Mp9@4736_d N_OUT8_Mp9@4736_g N_VDD_Mp9@4736_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4735 N_OUT9_Mn9@4735_d N_OUT8_Mn9@4735_g N_VSS_Mn9@4735_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4734 N_OUT9_Mn9@4734_d N_OUT8_Mn9@4734_g N_VSS_Mn9@4734_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4735 N_OUT9_Mp9@4735_d N_OUT8_Mp9@4735_g N_VDD_Mp9@4735_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4734 N_OUT9_Mp9@4734_d N_OUT8_Mp9@4734_g N_VDD_Mp9@4734_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4733 N_OUT9_Mn9@4733_d N_OUT8_Mn9@4733_g N_VSS_Mn9@4733_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4732 N_OUT9_Mn9@4732_d N_OUT8_Mn9@4732_g N_VSS_Mn9@4732_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4733 N_OUT9_Mp9@4733_d N_OUT8_Mp9@4733_g N_VDD_Mp9@4733_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4732 N_OUT9_Mp9@4732_d N_OUT8_Mp9@4732_g N_VDD_Mp9@4732_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4731 N_OUT9_Mn9@4731_d N_OUT8_Mn9@4731_g N_VSS_Mn9@4731_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4730 N_OUT9_Mn9@4730_d N_OUT8_Mn9@4730_g N_VSS_Mn9@4730_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4731 N_OUT9_Mp9@4731_d N_OUT8_Mp9@4731_g N_VDD_Mp9@4731_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4730 N_OUT9_Mp9@4730_d N_OUT8_Mp9@4730_g N_VDD_Mp9@4730_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4729 N_OUT9_Mn9@4729_d N_OUT8_Mn9@4729_g N_VSS_Mn9@4729_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4728 N_OUT9_Mn9@4728_d N_OUT8_Mn9@4728_g N_VSS_Mn9@4728_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4729 N_OUT9_Mp9@4729_d N_OUT8_Mp9@4729_g N_VDD_Mp9@4729_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4728 N_OUT9_Mp9@4728_d N_OUT8_Mp9@4728_g N_VDD_Mp9@4728_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4727 N_OUT9_Mn9@4727_d N_OUT8_Mn9@4727_g N_VSS_Mn9@4727_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4726 N_OUT9_Mn9@4726_d N_OUT8_Mn9@4726_g N_VSS_Mn9@4726_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4727 N_OUT9_Mp9@4727_d N_OUT8_Mp9@4727_g N_VDD_Mp9@4727_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4726 N_OUT9_Mp9@4726_d N_OUT8_Mp9@4726_g N_VDD_Mp9@4726_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4725 N_OUT9_Mn9@4725_d N_OUT8_Mn9@4725_g N_VSS_Mn9@4725_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4724 N_OUT9_Mn9@4724_d N_OUT8_Mn9@4724_g N_VSS_Mn9@4724_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4725 N_OUT9_Mp9@4725_d N_OUT8_Mp9@4725_g N_VDD_Mp9@4725_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4724 N_OUT9_Mp9@4724_d N_OUT8_Mp9@4724_g N_VDD_Mp9@4724_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4723 N_OUT9_Mn9@4723_d N_OUT8_Mn9@4723_g N_VSS_Mn9@4723_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4722 N_OUT9_Mn9@4722_d N_OUT8_Mn9@4722_g N_VSS_Mn9@4722_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4723 N_OUT9_Mp9@4723_d N_OUT8_Mp9@4723_g N_VDD_Mp9@4723_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4722 N_OUT9_Mp9@4722_d N_OUT8_Mp9@4722_g N_VDD_Mp9@4722_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4721 N_OUT9_Mn9@4721_d N_OUT8_Mn9@4721_g N_VSS_Mn9@4721_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4720 N_OUT9_Mn9@4720_d N_OUT8_Mn9@4720_g N_VSS_Mn9@4720_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4721 N_OUT9_Mp9@4721_d N_OUT8_Mp9@4721_g N_VDD_Mp9@4721_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4720 N_OUT9_Mp9@4720_d N_OUT8_Mp9@4720_g N_VDD_Mp9@4720_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4719 N_OUT9_Mn9@4719_d N_OUT8_Mn9@4719_g N_VSS_Mn9@4719_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4718 N_OUT9_Mn9@4718_d N_OUT8_Mn9@4718_g N_VSS_Mn9@4718_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4719 N_OUT9_Mp9@4719_d N_OUT8_Mp9@4719_g N_VDD_Mp9@4719_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4718 N_OUT9_Mp9@4718_d N_OUT8_Mp9@4718_g N_VDD_Mp9@4718_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4717 N_OUT9_Mn9@4717_d N_OUT8_Mn9@4717_g N_VSS_Mn9@4717_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4716 N_OUT9_Mn9@4716_d N_OUT8_Mn9@4716_g N_VSS_Mn9@4716_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4717 N_OUT9_Mp9@4717_d N_OUT8_Mp9@4717_g N_VDD_Mp9@4717_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4716 N_OUT9_Mp9@4716_d N_OUT8_Mp9@4716_g N_VDD_Mp9@4716_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4715 N_OUT9_Mn9@4715_d N_OUT8_Mn9@4715_g N_VSS_Mn9@4715_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4714 N_OUT9_Mn9@4714_d N_OUT8_Mn9@4714_g N_VSS_Mn9@4714_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4715 N_OUT9_Mp9@4715_d N_OUT8_Mp9@4715_g N_VDD_Mp9@4715_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4714 N_OUT9_Mp9@4714_d N_OUT8_Mp9@4714_g N_VDD_Mp9@4714_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4713 N_OUT9_Mn9@4713_d N_OUT8_Mn9@4713_g N_VSS_Mn9@4713_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4712 N_OUT9_Mn9@4712_d N_OUT8_Mn9@4712_g N_VSS_Mn9@4712_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4713 N_OUT9_Mp9@4713_d N_OUT8_Mp9@4713_g N_VDD_Mp9@4713_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4712 N_OUT9_Mp9@4712_d N_OUT8_Mp9@4712_g N_VDD_Mp9@4712_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4711 N_OUT9_Mn9@4711_d N_OUT8_Mn9@4711_g N_VSS_Mn9@4711_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4710 N_OUT9_Mn9@4710_d N_OUT8_Mn9@4710_g N_VSS_Mn9@4710_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4711 N_OUT9_Mp9@4711_d N_OUT8_Mp9@4711_g N_VDD_Mp9@4711_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4710 N_OUT9_Mp9@4710_d N_OUT8_Mp9@4710_g N_VDD_Mp9@4710_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4709 N_OUT9_Mn9@4709_d N_OUT8_Mn9@4709_g N_VSS_Mn9@4709_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4708 N_OUT9_Mn9@4708_d N_OUT8_Mn9@4708_g N_VSS_Mn9@4708_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4709 N_OUT9_Mp9@4709_d N_OUT8_Mp9@4709_g N_VDD_Mp9@4709_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4708 N_OUT9_Mp9@4708_d N_OUT8_Mp9@4708_g N_VDD_Mp9@4708_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4707 N_OUT9_Mn9@4707_d N_OUT8_Mn9@4707_g N_VSS_Mn9@4707_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4706 N_OUT9_Mn9@4706_d N_OUT8_Mn9@4706_g N_VSS_Mn9@4706_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4707 N_OUT9_Mp9@4707_d N_OUT8_Mp9@4707_g N_VDD_Mp9@4707_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4706 N_OUT9_Mp9@4706_d N_OUT8_Mp9@4706_g N_VDD_Mp9@4706_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4705 N_OUT9_Mn9@4705_d N_OUT8_Mn9@4705_g N_VSS_Mn9@4705_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4704 N_OUT9_Mn9@4704_d N_OUT8_Mn9@4704_g N_VSS_Mn9@4704_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4705 N_OUT9_Mp9@4705_d N_OUT8_Mp9@4705_g N_VDD_Mp9@4705_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4704 N_OUT9_Mp9@4704_d N_OUT8_Mp9@4704_g N_VDD_Mp9@4704_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4703 N_OUT9_Mn9@4703_d N_OUT8_Mn9@4703_g N_VSS_Mn9@4703_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4702 N_OUT9_Mn9@4702_d N_OUT8_Mn9@4702_g N_VSS_Mn9@4702_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4703 N_OUT9_Mp9@4703_d N_OUT8_Mp9@4703_g N_VDD_Mp9@4703_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4702 N_OUT9_Mp9@4702_d N_OUT8_Mp9@4702_g N_VDD_Mp9@4702_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4701 N_OUT9_Mn9@4701_d N_OUT8_Mn9@4701_g N_VSS_Mn9@4701_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4700 N_OUT9_Mn9@4700_d N_OUT8_Mn9@4700_g N_VSS_Mn9@4700_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4701 N_OUT9_Mp9@4701_d N_OUT8_Mp9@4701_g N_VDD_Mp9@4701_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4700 N_OUT9_Mp9@4700_d N_OUT8_Mp9@4700_g N_VDD_Mp9@4700_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4699 N_OUT9_Mn9@4699_d N_OUT8_Mn9@4699_g N_VSS_Mn9@4699_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4698 N_OUT9_Mn9@4698_d N_OUT8_Mn9@4698_g N_VSS_Mn9@4698_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4699 N_OUT9_Mp9@4699_d N_OUT8_Mp9@4699_g N_VDD_Mp9@4699_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4698 N_OUT9_Mp9@4698_d N_OUT8_Mp9@4698_g N_VDD_Mp9@4698_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4697 N_OUT9_Mn9@4697_d N_OUT8_Mn9@4697_g N_VSS_Mn9@4697_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4696 N_OUT9_Mn9@4696_d N_OUT8_Mn9@4696_g N_VSS_Mn9@4696_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4697 N_OUT9_Mp9@4697_d N_OUT8_Mp9@4697_g N_VDD_Mp9@4697_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4696 N_OUT9_Mp9@4696_d N_OUT8_Mp9@4696_g N_VDD_Mp9@4696_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4695 N_OUT9_Mn9@4695_d N_OUT8_Mn9@4695_g N_VSS_Mn9@4695_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4694 N_OUT9_Mn9@4694_d N_OUT8_Mn9@4694_g N_VSS_Mn9@4694_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4695 N_OUT9_Mp9@4695_d N_OUT8_Mp9@4695_g N_VDD_Mp9@4695_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4694 N_OUT9_Mp9@4694_d N_OUT8_Mp9@4694_g N_VDD_Mp9@4694_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4693 N_OUT9_Mn9@4693_d N_OUT8_Mn9@4693_g N_VSS_Mn9@4693_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4692 N_OUT9_Mn9@4692_d N_OUT8_Mn9@4692_g N_VSS_Mn9@4692_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4693 N_OUT9_Mp9@4693_d N_OUT8_Mp9@4693_g N_VDD_Mp9@4693_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4692 N_OUT9_Mp9@4692_d N_OUT8_Mp9@4692_g N_VDD_Mp9@4692_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4691 N_OUT9_Mn9@4691_d N_OUT8_Mn9@4691_g N_VSS_Mn9@4691_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4690 N_OUT9_Mn9@4690_d N_OUT8_Mn9@4690_g N_VSS_Mn9@4690_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4691 N_OUT9_Mp9@4691_d N_OUT8_Mp9@4691_g N_VDD_Mp9@4691_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4690 N_OUT9_Mp9@4690_d N_OUT8_Mp9@4690_g N_VDD_Mp9@4690_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4689 N_OUT9_Mn9@4689_d N_OUT8_Mn9@4689_g N_VSS_Mn9@4689_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4688 N_OUT9_Mn9@4688_d N_OUT8_Mn9@4688_g N_VSS_Mn9@4688_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4689 N_OUT9_Mp9@4689_d N_OUT8_Mp9@4689_g N_VDD_Mp9@4689_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4688 N_OUT9_Mp9@4688_d N_OUT8_Mp9@4688_g N_VDD_Mp9@4688_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4687 N_OUT9_Mn9@4687_d N_OUT8_Mn9@4687_g N_VSS_Mn9@4687_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4686 N_OUT9_Mn9@4686_d N_OUT8_Mn9@4686_g N_VSS_Mn9@4686_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4687 N_OUT9_Mp9@4687_d N_OUT8_Mp9@4687_g N_VDD_Mp9@4687_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4686 N_OUT9_Mp9@4686_d N_OUT8_Mp9@4686_g N_VDD_Mp9@4686_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4685 N_OUT9_Mn9@4685_d N_OUT8_Mn9@4685_g N_VSS_Mn9@4685_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4684 N_OUT9_Mn9@4684_d N_OUT8_Mn9@4684_g N_VSS_Mn9@4684_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4685 N_OUT9_Mp9@4685_d N_OUT8_Mp9@4685_g N_VDD_Mp9@4685_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4684 N_OUT9_Mp9@4684_d N_OUT8_Mp9@4684_g N_VDD_Mp9@4684_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4683 N_OUT9_Mn9@4683_d N_OUT8_Mn9@4683_g N_VSS_Mn9@4683_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4682 N_OUT9_Mn9@4682_d N_OUT8_Mn9@4682_g N_VSS_Mn9@4682_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4683 N_OUT9_Mp9@4683_d N_OUT8_Mp9@4683_g N_VDD_Mp9@4683_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4682 N_OUT9_Mp9@4682_d N_OUT8_Mp9@4682_g N_VDD_Mp9@4682_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4681 N_OUT9_Mn9@4681_d N_OUT8_Mn9@4681_g N_VSS_Mn9@4681_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4680 N_OUT9_Mn9@4680_d N_OUT8_Mn9@4680_g N_VSS_Mn9@4680_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4681 N_OUT9_Mp9@4681_d N_OUT8_Mp9@4681_g N_VDD_Mp9@4681_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4680 N_OUT9_Mp9@4680_d N_OUT8_Mp9@4680_g N_VDD_Mp9@4680_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4679 N_OUT9_Mn9@4679_d N_OUT8_Mn9@4679_g N_VSS_Mn9@4679_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4678 N_OUT9_Mn9@4678_d N_OUT8_Mn9@4678_g N_VSS_Mn9@4678_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4679 N_OUT9_Mp9@4679_d N_OUT8_Mp9@4679_g N_VDD_Mp9@4679_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4678 N_OUT9_Mp9@4678_d N_OUT8_Mp9@4678_g N_VDD_Mp9@4678_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4677 N_OUT9_Mn9@4677_d N_OUT8_Mn9@4677_g N_VSS_Mn9@4677_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4676 N_OUT9_Mn9@4676_d N_OUT8_Mn9@4676_g N_VSS_Mn9@4676_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4677 N_OUT9_Mp9@4677_d N_OUT8_Mp9@4677_g N_VDD_Mp9@4677_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4676 N_OUT9_Mp9@4676_d N_OUT8_Mp9@4676_g N_VDD_Mp9@4676_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4675 N_OUT9_Mn9@4675_d N_OUT8_Mn9@4675_g N_VSS_Mn9@4675_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4674 N_OUT9_Mn9@4674_d N_OUT8_Mn9@4674_g N_VSS_Mn9@4674_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4675 N_OUT9_Mp9@4675_d N_OUT8_Mp9@4675_g N_VDD_Mp9@4675_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4674 N_OUT9_Mp9@4674_d N_OUT8_Mp9@4674_g N_VDD_Mp9@4674_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4673 N_OUT9_Mn9@4673_d N_OUT8_Mn9@4673_g N_VSS_Mn9@4673_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4672 N_OUT9_Mn9@4672_d N_OUT8_Mn9@4672_g N_VSS_Mn9@4672_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4673 N_OUT9_Mp9@4673_d N_OUT8_Mp9@4673_g N_VDD_Mp9@4673_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4672 N_OUT9_Mp9@4672_d N_OUT8_Mp9@4672_g N_VDD_Mp9@4672_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4671 N_OUT9_Mn9@4671_d N_OUT8_Mn9@4671_g N_VSS_Mn9@4671_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4670 N_OUT9_Mn9@4670_d N_OUT8_Mn9@4670_g N_VSS_Mn9@4670_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4671 N_OUT9_Mp9@4671_d N_OUT8_Mp9@4671_g N_VDD_Mp9@4671_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4670 N_OUT9_Mp9@4670_d N_OUT8_Mp9@4670_g N_VDD_Mp9@4670_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4669 N_OUT9_Mn9@4669_d N_OUT8_Mn9@4669_g N_VSS_Mn9@4669_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4668 N_OUT9_Mn9@4668_d N_OUT8_Mn9@4668_g N_VSS_Mn9@4668_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4669 N_OUT9_Mp9@4669_d N_OUT8_Mp9@4669_g N_VDD_Mp9@4669_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4668 N_OUT9_Mp9@4668_d N_OUT8_Mp9@4668_g N_VDD_Mp9@4668_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4667 N_OUT9_Mn9@4667_d N_OUT8_Mn9@4667_g N_VSS_Mn9@4667_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4666 N_OUT9_Mn9@4666_d N_OUT8_Mn9@4666_g N_VSS_Mn9@4666_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4667 N_OUT9_Mp9@4667_d N_OUT8_Mp9@4667_g N_VDD_Mp9@4667_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4666 N_OUT9_Mp9@4666_d N_OUT8_Mp9@4666_g N_VDD_Mp9@4666_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4665 N_OUT9_Mn9@4665_d N_OUT8_Mn9@4665_g N_VSS_Mn9@4665_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4664 N_OUT9_Mn9@4664_d N_OUT8_Mn9@4664_g N_VSS_Mn9@4664_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4665 N_OUT9_Mp9@4665_d N_OUT8_Mp9@4665_g N_VDD_Mp9@4665_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4664 N_OUT9_Mp9@4664_d N_OUT8_Mp9@4664_g N_VDD_Mp9@4664_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4663 N_OUT9_Mn9@4663_d N_OUT8_Mn9@4663_g N_VSS_Mn9@4663_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4662 N_OUT9_Mn9@4662_d N_OUT8_Mn9@4662_g N_VSS_Mn9@4662_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4663 N_OUT9_Mp9@4663_d N_OUT8_Mp9@4663_g N_VDD_Mp9@4663_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4662 N_OUT9_Mp9@4662_d N_OUT8_Mp9@4662_g N_VDD_Mp9@4662_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4661 N_OUT9_Mn9@4661_d N_OUT8_Mn9@4661_g N_VSS_Mn9@4661_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4660 N_OUT9_Mn9@4660_d N_OUT8_Mn9@4660_g N_VSS_Mn9@4660_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4661 N_OUT9_Mp9@4661_d N_OUT8_Mp9@4661_g N_VDD_Mp9@4661_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4660 N_OUT9_Mp9@4660_d N_OUT8_Mp9@4660_g N_VDD_Mp9@4660_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4659 N_OUT9_Mn9@4659_d N_OUT8_Mn9@4659_g N_VSS_Mn9@4659_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4658 N_OUT9_Mn9@4658_d N_OUT8_Mn9@4658_g N_VSS_Mn9@4658_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4659 N_OUT9_Mp9@4659_d N_OUT8_Mp9@4659_g N_VDD_Mp9@4659_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4658 N_OUT9_Mp9@4658_d N_OUT8_Mp9@4658_g N_VDD_Mp9@4658_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4657 N_OUT9_Mn9@4657_d N_OUT8_Mn9@4657_g N_VSS_Mn9@4657_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4656 N_OUT9_Mn9@4656_d N_OUT8_Mn9@4656_g N_VSS_Mn9@4656_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4657 N_OUT9_Mp9@4657_d N_OUT8_Mp9@4657_g N_VDD_Mp9@4657_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4656 N_OUT9_Mp9@4656_d N_OUT8_Mp9@4656_g N_VDD_Mp9@4656_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4655 N_OUT9_Mn9@4655_d N_OUT8_Mn9@4655_g N_VSS_Mn9@4655_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4654 N_OUT9_Mn9@4654_d N_OUT8_Mn9@4654_g N_VSS_Mn9@4654_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4655 N_OUT9_Mp9@4655_d N_OUT8_Mp9@4655_g N_VDD_Mp9@4655_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4654 N_OUT9_Mp9@4654_d N_OUT8_Mp9@4654_g N_VDD_Mp9@4654_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4653 N_OUT9_Mn9@4653_d N_OUT8_Mn9@4653_g N_VSS_Mn9@4653_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4652 N_OUT9_Mn9@4652_d N_OUT8_Mn9@4652_g N_VSS_Mn9@4652_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4653 N_OUT9_Mp9@4653_d N_OUT8_Mp9@4653_g N_VDD_Mp9@4653_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4652 N_OUT9_Mp9@4652_d N_OUT8_Mp9@4652_g N_VDD_Mp9@4652_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4651 N_OUT9_Mn9@4651_d N_OUT8_Mn9@4651_g N_VSS_Mn9@4651_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4650 N_OUT9_Mn9@4650_d N_OUT8_Mn9@4650_g N_VSS_Mn9@4650_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4651 N_OUT9_Mp9@4651_d N_OUT8_Mp9@4651_g N_VDD_Mp9@4651_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4650 N_OUT9_Mp9@4650_d N_OUT8_Mp9@4650_g N_VDD_Mp9@4650_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4649 N_OUT9_Mn9@4649_d N_OUT8_Mn9@4649_g N_VSS_Mn9@4649_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4648 N_OUT9_Mn9@4648_d N_OUT8_Mn9@4648_g N_VSS_Mn9@4648_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4649 N_OUT9_Mp9@4649_d N_OUT8_Mp9@4649_g N_VDD_Mp9@4649_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4648 N_OUT9_Mp9@4648_d N_OUT8_Mp9@4648_g N_VDD_Mp9@4648_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4647 N_OUT9_Mn9@4647_d N_OUT8_Mn9@4647_g N_VSS_Mn9@4647_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4646 N_OUT9_Mn9@4646_d N_OUT8_Mn9@4646_g N_VSS_Mn9@4646_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4647 N_OUT9_Mp9@4647_d N_OUT8_Mp9@4647_g N_VDD_Mp9@4647_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4646 N_OUT9_Mp9@4646_d N_OUT8_Mp9@4646_g N_VDD_Mp9@4646_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4645 N_OUT9_Mn9@4645_d N_OUT8_Mn9@4645_g N_VSS_Mn9@4645_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4644 N_OUT9_Mn9@4644_d N_OUT8_Mn9@4644_g N_VSS_Mn9@4644_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4645 N_OUT9_Mp9@4645_d N_OUT8_Mp9@4645_g N_VDD_Mp9@4645_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4644 N_OUT9_Mp9@4644_d N_OUT8_Mp9@4644_g N_VDD_Mp9@4644_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4643 N_OUT9_Mn9@4643_d N_OUT8_Mn9@4643_g N_VSS_Mn9@4643_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4642 N_OUT9_Mn9@4642_d N_OUT8_Mn9@4642_g N_VSS_Mn9@4642_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4643 N_OUT9_Mp9@4643_d N_OUT8_Mp9@4643_g N_VDD_Mp9@4643_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4642 N_OUT9_Mp9@4642_d N_OUT8_Mp9@4642_g N_VDD_Mp9@4642_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4641 N_OUT9_Mn9@4641_d N_OUT8_Mn9@4641_g N_VSS_Mn9@4641_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4640 N_OUT9_Mn9@4640_d N_OUT8_Mn9@4640_g N_VSS_Mn9@4640_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4641 N_OUT9_Mp9@4641_d N_OUT8_Mp9@4641_g N_VDD_Mp9@4641_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4640 N_OUT9_Mp9@4640_d N_OUT8_Mp9@4640_g N_VDD_Mp9@4640_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4639 N_OUT9_Mn9@4639_d N_OUT8_Mn9@4639_g N_VSS_Mn9@4639_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4638 N_OUT9_Mn9@4638_d N_OUT8_Mn9@4638_g N_VSS_Mn9@4638_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4639 N_OUT9_Mp9@4639_d N_OUT8_Mp9@4639_g N_VDD_Mp9@4639_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4638 N_OUT9_Mp9@4638_d N_OUT8_Mp9@4638_g N_VDD_Mp9@4638_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4637 N_OUT9_Mn9@4637_d N_OUT8_Mn9@4637_g N_VSS_Mn9@4637_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4636 N_OUT9_Mn9@4636_d N_OUT8_Mn9@4636_g N_VSS_Mn9@4636_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4637 N_OUT9_Mp9@4637_d N_OUT8_Mp9@4637_g N_VDD_Mp9@4637_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4636 N_OUT9_Mp9@4636_d N_OUT8_Mp9@4636_g N_VDD_Mp9@4636_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4635 N_OUT9_Mn9@4635_d N_OUT8_Mn9@4635_g N_VSS_Mn9@4635_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4634 N_OUT9_Mn9@4634_d N_OUT8_Mn9@4634_g N_VSS_Mn9@4634_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4635 N_OUT9_Mp9@4635_d N_OUT8_Mp9@4635_g N_VDD_Mp9@4635_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4634 N_OUT9_Mp9@4634_d N_OUT8_Mp9@4634_g N_VDD_Mp9@4634_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4633 N_OUT9_Mn9@4633_d N_OUT8_Mn9@4633_g N_VSS_Mn9@4633_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4632 N_OUT9_Mn9@4632_d N_OUT8_Mn9@4632_g N_VSS_Mn9@4632_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4633 N_OUT9_Mp9@4633_d N_OUT8_Mp9@4633_g N_VDD_Mp9@4633_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4632 N_OUT9_Mp9@4632_d N_OUT8_Mp9@4632_g N_VDD_Mp9@4632_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4631 N_OUT9_Mn9@4631_d N_OUT8_Mn9@4631_g N_VSS_Mn9@4631_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4630 N_OUT9_Mn9@4630_d N_OUT8_Mn9@4630_g N_VSS_Mn9@4630_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4631 N_OUT9_Mp9@4631_d N_OUT8_Mp9@4631_g N_VDD_Mp9@4631_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4630 N_OUT9_Mp9@4630_d N_OUT8_Mp9@4630_g N_VDD_Mp9@4630_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4629 N_OUT9_Mn9@4629_d N_OUT8_Mn9@4629_g N_VSS_Mn9@4629_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4628 N_OUT9_Mn9@4628_d N_OUT8_Mn9@4628_g N_VSS_Mn9@4628_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4629 N_OUT9_Mp9@4629_d N_OUT8_Mp9@4629_g N_VDD_Mp9@4629_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4628 N_OUT9_Mp9@4628_d N_OUT8_Mp9@4628_g N_VDD_Mp9@4628_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4627 N_OUT9_Mn9@4627_d N_OUT8_Mn9@4627_g N_VSS_Mn9@4627_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4626 N_OUT9_Mn9@4626_d N_OUT8_Mn9@4626_g N_VSS_Mn9@4626_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4627 N_OUT9_Mp9@4627_d N_OUT8_Mp9@4627_g N_VDD_Mp9@4627_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4626 N_OUT9_Mp9@4626_d N_OUT8_Mp9@4626_g N_VDD_Mp9@4626_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4625 N_OUT9_Mn9@4625_d N_OUT8_Mn9@4625_g N_VSS_Mn9@4625_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4624 N_OUT9_Mn9@4624_d N_OUT8_Mn9@4624_g N_VSS_Mn9@4624_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4625 N_OUT9_Mp9@4625_d N_OUT8_Mp9@4625_g N_VDD_Mp9@4625_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4624 N_OUT9_Mp9@4624_d N_OUT8_Mp9@4624_g N_VDD_Mp9@4624_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4623 N_OUT9_Mn9@4623_d N_OUT8_Mn9@4623_g N_VSS_Mn9@4623_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4622 N_OUT9_Mn9@4622_d N_OUT8_Mn9@4622_g N_VSS_Mn9@4622_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4623 N_OUT9_Mp9@4623_d N_OUT8_Mp9@4623_g N_VDD_Mp9@4623_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4622 N_OUT9_Mp9@4622_d N_OUT8_Mp9@4622_g N_VDD_Mp9@4622_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4621 N_OUT9_Mn9@4621_d N_OUT8_Mn9@4621_g N_VSS_Mn9@4621_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4620 N_OUT9_Mn9@4620_d N_OUT8_Mn9@4620_g N_VSS_Mn9@4620_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4621 N_OUT9_Mp9@4621_d N_OUT8_Mp9@4621_g N_VDD_Mp9@4621_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4620 N_OUT9_Mp9@4620_d N_OUT8_Mp9@4620_g N_VDD_Mp9@4620_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4619 N_OUT9_Mn9@4619_d N_OUT8_Mn9@4619_g N_VSS_Mn9@4619_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4618 N_OUT9_Mn9@4618_d N_OUT8_Mn9@4618_g N_VSS_Mn9@4618_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4619 N_OUT9_Mp9@4619_d N_OUT8_Mp9@4619_g N_VDD_Mp9@4619_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4618 N_OUT9_Mp9@4618_d N_OUT8_Mp9@4618_g N_VDD_Mp9@4618_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4617 N_OUT9_Mn9@4617_d N_OUT8_Mn9@4617_g N_VSS_Mn9@4617_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4616 N_OUT9_Mn9@4616_d N_OUT8_Mn9@4616_g N_VSS_Mn9@4616_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4617 N_OUT9_Mp9@4617_d N_OUT8_Mp9@4617_g N_VDD_Mp9@4617_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4616 N_OUT9_Mp9@4616_d N_OUT8_Mp9@4616_g N_VDD_Mp9@4616_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4615 N_OUT9_Mn9@4615_d N_OUT8_Mn9@4615_g N_VSS_Mn9@4615_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4614 N_OUT9_Mn9@4614_d N_OUT8_Mn9@4614_g N_VSS_Mn9@4614_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4615 N_OUT9_Mp9@4615_d N_OUT8_Mp9@4615_g N_VDD_Mp9@4615_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4614 N_OUT9_Mp9@4614_d N_OUT8_Mp9@4614_g N_VDD_Mp9@4614_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4613 N_OUT9_Mn9@4613_d N_OUT8_Mn9@4613_g N_VSS_Mn9@4613_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4612 N_OUT9_Mn9@4612_d N_OUT8_Mn9@4612_g N_VSS_Mn9@4612_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4613 N_OUT9_Mp9@4613_d N_OUT8_Mp9@4613_g N_VDD_Mp9@4613_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4612 N_OUT9_Mp9@4612_d N_OUT8_Mp9@4612_g N_VDD_Mp9@4612_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4611 N_OUT9_Mn9@4611_d N_OUT8_Mn9@4611_g N_VSS_Mn9@4611_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4610 N_OUT9_Mn9@4610_d N_OUT8_Mn9@4610_g N_VSS_Mn9@4610_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4611 N_OUT9_Mp9@4611_d N_OUT8_Mp9@4611_g N_VDD_Mp9@4611_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4610 N_OUT9_Mp9@4610_d N_OUT8_Mp9@4610_g N_VDD_Mp9@4610_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3585 N_OUT8_Mn8@3585_d N_OUT7_Mn8@3585_g N_VSS_Mn8@3585_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3584 N_OUT8_Mn8@3584_d N_OUT7_Mn8@3584_g N_VSS_Mn8@3584_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3585 N_OUT8_Mp8@3585_d N_OUT7_Mp8@3585_g N_VDD_Mp8@3585_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3584 N_OUT8_Mp8@3584_d N_OUT7_Mp8@3584_g N_VDD_Mp8@3584_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3583 N_OUT8_Mn8@3583_d N_OUT7_Mn8@3583_g N_VSS_Mn8@3583_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3582 N_OUT8_Mn8@3582_d N_OUT7_Mn8@3582_g N_VSS_Mn8@3582_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3583 N_OUT8_Mp8@3583_d N_OUT7_Mp8@3583_g N_VDD_Mp8@3583_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3582 N_OUT8_Mp8@3582_d N_OUT7_Mp8@3582_g N_VDD_Mp8@3582_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3581 N_OUT8_Mn8@3581_d N_OUT7_Mn8@3581_g N_VSS_Mn8@3581_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3580 N_OUT8_Mn8@3580_d N_OUT7_Mn8@3580_g N_VSS_Mn8@3580_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3581 N_OUT8_Mp8@3581_d N_OUT7_Mp8@3581_g N_VDD_Mp8@3581_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3580 N_OUT8_Mp8@3580_d N_OUT7_Mp8@3580_g N_VDD_Mp8@3580_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3579 N_OUT8_Mn8@3579_d N_OUT7_Mn8@3579_g N_VSS_Mn8@3579_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3578 N_OUT8_Mn8@3578_d N_OUT7_Mn8@3578_g N_VSS_Mn8@3578_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3579 N_OUT8_Mp8@3579_d N_OUT7_Mp8@3579_g N_VDD_Mp8@3579_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3578 N_OUT8_Mp8@3578_d N_OUT7_Mp8@3578_g N_VDD_Mp8@3578_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3577 N_OUT8_Mn8@3577_d N_OUT7_Mn8@3577_g N_VSS_Mn8@3577_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3576 N_OUT8_Mn8@3576_d N_OUT7_Mn8@3576_g N_VSS_Mn8@3576_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3577 N_OUT8_Mp8@3577_d N_OUT7_Mp8@3577_g N_VDD_Mp8@3577_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3576 N_OUT8_Mp8@3576_d N_OUT7_Mp8@3576_g N_VDD_Mp8@3576_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3575 N_OUT8_Mn8@3575_d N_OUT7_Mn8@3575_g N_VSS_Mn8@3575_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3574 N_OUT8_Mn8@3574_d N_OUT7_Mn8@3574_g N_VSS_Mn8@3574_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3575 N_OUT8_Mp8@3575_d N_OUT7_Mp8@3575_g N_VDD_Mp8@3575_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3574 N_OUT8_Mp8@3574_d N_OUT7_Mp8@3574_g N_VDD_Mp8@3574_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3573 N_OUT8_Mn8@3573_d N_OUT7_Mn8@3573_g N_VSS_Mn8@3573_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3572 N_OUT8_Mn8@3572_d N_OUT7_Mn8@3572_g N_VSS_Mn8@3572_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3573 N_OUT8_Mp8@3573_d N_OUT7_Mp8@3573_g N_VDD_Mp8@3573_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3572 N_OUT8_Mp8@3572_d N_OUT7_Mp8@3572_g N_VDD_Mp8@3572_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3571 N_OUT8_Mn8@3571_d N_OUT7_Mn8@3571_g N_VSS_Mn8@3571_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3570 N_OUT8_Mn8@3570_d N_OUT7_Mn8@3570_g N_VSS_Mn8@3570_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3571 N_OUT8_Mp8@3571_d N_OUT7_Mp8@3571_g N_VDD_Mp8@3571_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3570 N_OUT8_Mp8@3570_d N_OUT7_Mp8@3570_g N_VDD_Mp8@3570_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3569 N_OUT8_Mn8@3569_d N_OUT7_Mn8@3569_g N_VSS_Mn8@3569_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3568 N_OUT8_Mn8@3568_d N_OUT7_Mn8@3568_g N_VSS_Mn8@3568_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3569 N_OUT8_Mp8@3569_d N_OUT7_Mp8@3569_g N_VDD_Mp8@3569_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3568 N_OUT8_Mp8@3568_d N_OUT7_Mp8@3568_g N_VDD_Mp8@3568_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3567 N_OUT8_Mn8@3567_d N_OUT7_Mn8@3567_g N_VSS_Mn8@3567_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3566 N_OUT8_Mn8@3566_d N_OUT7_Mn8@3566_g N_VSS_Mn8@3566_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3567 N_OUT8_Mp8@3567_d N_OUT7_Mp8@3567_g N_VDD_Mp8@3567_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3566 N_OUT8_Mp8@3566_d N_OUT7_Mp8@3566_g N_VDD_Mp8@3566_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3565 N_OUT8_Mn8@3565_d N_OUT7_Mn8@3565_g N_VSS_Mn8@3565_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3564 N_OUT8_Mn8@3564_d N_OUT7_Mn8@3564_g N_VSS_Mn8@3564_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3565 N_OUT8_Mp8@3565_d N_OUT7_Mp8@3565_g N_VDD_Mp8@3565_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3564 N_OUT8_Mp8@3564_d N_OUT7_Mp8@3564_g N_VDD_Mp8@3564_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3563 N_OUT8_Mn8@3563_d N_OUT7_Mn8@3563_g N_VSS_Mn8@3563_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3562 N_OUT8_Mn8@3562_d N_OUT7_Mn8@3562_g N_VSS_Mn8@3562_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3563 N_OUT8_Mp8@3563_d N_OUT7_Mp8@3563_g N_VDD_Mp8@3563_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3562 N_OUT8_Mp8@3562_d N_OUT7_Mp8@3562_g N_VDD_Mp8@3562_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3561 N_OUT8_Mn8@3561_d N_OUT7_Mn8@3561_g N_VSS_Mn8@3561_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3560 N_OUT8_Mn8@3560_d N_OUT7_Mn8@3560_g N_VSS_Mn8@3560_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3561 N_OUT8_Mp8@3561_d N_OUT7_Mp8@3561_g N_VDD_Mp8@3561_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3560 N_OUT8_Mp8@3560_d N_OUT7_Mp8@3560_g N_VDD_Mp8@3560_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3559 N_OUT8_Mn8@3559_d N_OUT7_Mn8@3559_g N_VSS_Mn8@3559_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3558 N_OUT8_Mn8@3558_d N_OUT7_Mn8@3558_g N_VSS_Mn8@3558_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3559 N_OUT8_Mp8@3559_d N_OUT7_Mp8@3559_g N_VDD_Mp8@3559_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3558 N_OUT8_Mp8@3558_d N_OUT7_Mp8@3558_g N_VDD_Mp8@3558_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3557 N_OUT8_Mn8@3557_d N_OUT7_Mn8@3557_g N_VSS_Mn8@3557_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3556 N_OUT8_Mn8@3556_d N_OUT7_Mn8@3556_g N_VSS_Mn8@3556_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3557 N_OUT8_Mp8@3557_d N_OUT7_Mp8@3557_g N_VDD_Mp8@3557_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3556 N_OUT8_Mp8@3556_d N_OUT7_Mp8@3556_g N_VDD_Mp8@3556_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3555 N_OUT8_Mn8@3555_d N_OUT7_Mn8@3555_g N_VSS_Mn8@3555_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3554 N_OUT8_Mn8@3554_d N_OUT7_Mn8@3554_g N_VSS_Mn8@3554_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3555 N_OUT8_Mp8@3555_d N_OUT7_Mp8@3555_g N_VDD_Mp8@3555_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3554 N_OUT8_Mp8@3554_d N_OUT7_Mp8@3554_g N_VDD_Mp8@3554_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3553 N_OUT8_Mn8@3553_d N_OUT7_Mn8@3553_g N_VSS_Mn8@3553_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3552 N_OUT8_Mn8@3552_d N_OUT7_Mn8@3552_g N_VSS_Mn8@3552_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3553 N_OUT8_Mp8@3553_d N_OUT7_Mp8@3553_g N_VDD_Mp8@3553_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3552 N_OUT8_Mp8@3552_d N_OUT7_Mp8@3552_g N_VDD_Mp8@3552_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3551 N_OUT8_Mn8@3551_d N_OUT7_Mn8@3551_g N_VSS_Mn8@3551_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3550 N_OUT8_Mn8@3550_d N_OUT7_Mn8@3550_g N_VSS_Mn8@3550_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3551 N_OUT8_Mp8@3551_d N_OUT7_Mp8@3551_g N_VDD_Mp8@3551_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3550 N_OUT8_Mp8@3550_d N_OUT7_Mp8@3550_g N_VDD_Mp8@3550_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3549 N_OUT8_Mn8@3549_d N_OUT7_Mn8@3549_g N_VSS_Mn8@3549_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3548 N_OUT8_Mn8@3548_d N_OUT7_Mn8@3548_g N_VSS_Mn8@3548_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3549 N_OUT8_Mp8@3549_d N_OUT7_Mp8@3549_g N_VDD_Mp8@3549_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3548 N_OUT8_Mp8@3548_d N_OUT7_Mp8@3548_g N_VDD_Mp8@3548_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3547 N_OUT8_Mn8@3547_d N_OUT7_Mn8@3547_g N_VSS_Mn8@3547_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3546 N_OUT8_Mn8@3546_d N_OUT7_Mn8@3546_g N_VSS_Mn8@3546_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3547 N_OUT8_Mp8@3547_d N_OUT7_Mp8@3547_g N_VDD_Mp8@3547_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3546 N_OUT8_Mp8@3546_d N_OUT7_Mp8@3546_g N_VDD_Mp8@3546_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3545 N_OUT8_Mn8@3545_d N_OUT7_Mn8@3545_g N_VSS_Mn8@3545_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3544 N_OUT8_Mn8@3544_d N_OUT7_Mn8@3544_g N_VSS_Mn8@3544_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3545 N_OUT8_Mp8@3545_d N_OUT7_Mp8@3545_g N_VDD_Mp8@3545_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3544 N_OUT8_Mp8@3544_d N_OUT7_Mp8@3544_g N_VDD_Mp8@3544_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3543 N_OUT8_Mn8@3543_d N_OUT7_Mn8@3543_g N_VSS_Mn8@3543_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3542 N_OUT8_Mn8@3542_d N_OUT7_Mn8@3542_g N_VSS_Mn8@3542_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3543 N_OUT8_Mp8@3543_d N_OUT7_Mp8@3543_g N_VDD_Mp8@3543_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3542 N_OUT8_Mp8@3542_d N_OUT7_Mp8@3542_g N_VDD_Mp8@3542_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3541 N_OUT8_Mn8@3541_d N_OUT7_Mn8@3541_g N_VSS_Mn8@3541_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3540 N_OUT8_Mn8@3540_d N_OUT7_Mn8@3540_g N_VSS_Mn8@3540_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3541 N_OUT8_Mp8@3541_d N_OUT7_Mp8@3541_g N_VDD_Mp8@3541_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3540 N_OUT8_Mp8@3540_d N_OUT7_Mp8@3540_g N_VDD_Mp8@3540_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3539 N_OUT8_Mn8@3539_d N_OUT7_Mn8@3539_g N_VSS_Mn8@3539_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3538 N_OUT8_Mn8@3538_d N_OUT7_Mn8@3538_g N_VSS_Mn8@3538_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3539 N_OUT8_Mp8@3539_d N_OUT7_Mp8@3539_g N_VDD_Mp8@3539_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3538 N_OUT8_Mp8@3538_d N_OUT7_Mp8@3538_g N_VDD_Mp8@3538_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3537 N_OUT8_Mn8@3537_d N_OUT7_Mn8@3537_g N_VSS_Mn8@3537_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3536 N_OUT8_Mn8@3536_d N_OUT7_Mn8@3536_g N_VSS_Mn8@3536_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3537 N_OUT8_Mp8@3537_d N_OUT7_Mp8@3537_g N_VDD_Mp8@3537_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3536 N_OUT8_Mp8@3536_d N_OUT7_Mp8@3536_g N_VDD_Mp8@3536_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3535 N_OUT8_Mn8@3535_d N_OUT7_Mn8@3535_g N_VSS_Mn8@3535_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3534 N_OUT8_Mn8@3534_d N_OUT7_Mn8@3534_g N_VSS_Mn8@3534_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3535 N_OUT8_Mp8@3535_d N_OUT7_Mp8@3535_g N_VDD_Mp8@3535_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3534 N_OUT8_Mp8@3534_d N_OUT7_Mp8@3534_g N_VDD_Mp8@3534_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3533 N_OUT8_Mn8@3533_d N_OUT7_Mn8@3533_g N_VSS_Mn8@3533_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3532 N_OUT8_Mn8@3532_d N_OUT7_Mn8@3532_g N_VSS_Mn8@3532_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3533 N_OUT8_Mp8@3533_d N_OUT7_Mp8@3533_g N_VDD_Mp8@3533_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3532 N_OUT8_Mp8@3532_d N_OUT7_Mp8@3532_g N_VDD_Mp8@3532_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3531 N_OUT8_Mn8@3531_d N_OUT7_Mn8@3531_g N_VSS_Mn8@3531_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3530 N_OUT8_Mn8@3530_d N_OUT7_Mn8@3530_g N_VSS_Mn8@3530_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3531 N_OUT8_Mp8@3531_d N_OUT7_Mp8@3531_g N_VDD_Mp8@3531_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3530 N_OUT8_Mp8@3530_d N_OUT7_Mp8@3530_g N_VDD_Mp8@3530_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3529 N_OUT8_Mn8@3529_d N_OUT7_Mn8@3529_g N_VSS_Mn8@3529_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3528 N_OUT8_Mn8@3528_d N_OUT7_Mn8@3528_g N_VSS_Mn8@3528_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3529 N_OUT8_Mp8@3529_d N_OUT7_Mp8@3529_g N_VDD_Mp8@3529_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3528 N_OUT8_Mp8@3528_d N_OUT7_Mp8@3528_g N_VDD_Mp8@3528_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3527 N_OUT8_Mn8@3527_d N_OUT7_Mn8@3527_g N_VSS_Mn8@3527_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3526 N_OUT8_Mn8@3526_d N_OUT7_Mn8@3526_g N_VSS_Mn8@3526_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3527 N_OUT8_Mp8@3527_d N_OUT7_Mp8@3527_g N_VDD_Mp8@3527_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3526 N_OUT8_Mp8@3526_d N_OUT7_Mp8@3526_g N_VDD_Mp8@3526_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3525 N_OUT8_Mn8@3525_d N_OUT7_Mn8@3525_g N_VSS_Mn8@3525_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3524 N_OUT8_Mn8@3524_d N_OUT7_Mn8@3524_g N_VSS_Mn8@3524_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3525 N_OUT8_Mp8@3525_d N_OUT7_Mp8@3525_g N_VDD_Mp8@3525_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3524 N_OUT8_Mp8@3524_d N_OUT7_Mp8@3524_g N_VDD_Mp8@3524_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3523 N_OUT8_Mn8@3523_d N_OUT7_Mn8@3523_g N_VSS_Mn8@3523_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3522 N_OUT8_Mn8@3522_d N_OUT7_Mn8@3522_g N_VSS_Mn8@3522_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3523 N_OUT8_Mp8@3523_d N_OUT7_Mp8@3523_g N_VDD_Mp8@3523_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3522 N_OUT8_Mp8@3522_d N_OUT7_Mp8@3522_g N_VDD_Mp8@3522_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3521 N_OUT8_Mn8@3521_d N_OUT7_Mn8@3521_g N_VSS_Mn8@3521_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3520 N_OUT8_Mn8@3520_d N_OUT7_Mn8@3520_g N_VSS_Mn8@3520_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3521 N_OUT8_Mp8@3521_d N_OUT7_Mp8@3521_g N_VDD_Mp8@3521_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3520 N_OUT8_Mp8@3520_d N_OUT7_Mp8@3520_g N_VDD_Mp8@3520_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3519 N_OUT8_Mn8@3519_d N_OUT7_Mn8@3519_g N_VSS_Mn8@3519_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3518 N_OUT8_Mn8@3518_d N_OUT7_Mn8@3518_g N_VSS_Mn8@3518_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3519 N_OUT8_Mp8@3519_d N_OUT7_Mp8@3519_g N_VDD_Mp8@3519_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3518 N_OUT8_Mp8@3518_d N_OUT7_Mp8@3518_g N_VDD_Mp8@3518_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3517 N_OUT8_Mn8@3517_d N_OUT7_Mn8@3517_g N_VSS_Mn8@3517_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3516 N_OUT8_Mn8@3516_d N_OUT7_Mn8@3516_g N_VSS_Mn8@3516_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3517 N_OUT8_Mp8@3517_d N_OUT7_Mp8@3517_g N_VDD_Mp8@3517_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3516 N_OUT8_Mp8@3516_d N_OUT7_Mp8@3516_g N_VDD_Mp8@3516_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3515 N_OUT8_Mn8@3515_d N_OUT7_Mn8@3515_g N_VSS_Mn8@3515_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3514 N_OUT8_Mn8@3514_d N_OUT7_Mn8@3514_g N_VSS_Mn8@3514_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3515 N_OUT8_Mp8@3515_d N_OUT7_Mp8@3515_g N_VDD_Mp8@3515_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3514 N_OUT8_Mp8@3514_d N_OUT7_Mp8@3514_g N_VDD_Mp8@3514_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3513 N_OUT8_Mn8@3513_d N_OUT7_Mn8@3513_g N_VSS_Mn8@3513_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3512 N_OUT8_Mn8@3512_d N_OUT7_Mn8@3512_g N_VSS_Mn8@3512_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3513 N_OUT8_Mp8@3513_d N_OUT7_Mp8@3513_g N_VDD_Mp8@3513_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3512 N_OUT8_Mp8@3512_d N_OUT7_Mp8@3512_g N_VDD_Mp8@3512_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3511 N_OUT8_Mn8@3511_d N_OUT7_Mn8@3511_g N_VSS_Mn8@3511_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3510 N_OUT8_Mn8@3510_d N_OUT7_Mn8@3510_g N_VSS_Mn8@3510_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3511 N_OUT8_Mp8@3511_d N_OUT7_Mp8@3511_g N_VDD_Mp8@3511_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3510 N_OUT8_Mp8@3510_d N_OUT7_Mp8@3510_g N_VDD_Mp8@3510_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3509 N_OUT8_Mn8@3509_d N_OUT7_Mn8@3509_g N_VSS_Mn8@3509_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3508 N_OUT8_Mn8@3508_d N_OUT7_Mn8@3508_g N_VSS_Mn8@3508_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3509 N_OUT8_Mp8@3509_d N_OUT7_Mp8@3509_g N_VDD_Mp8@3509_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3508 N_OUT8_Mp8@3508_d N_OUT7_Mp8@3508_g N_VDD_Mp8@3508_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3507 N_OUT8_Mn8@3507_d N_OUT7_Mn8@3507_g N_VSS_Mn8@3507_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3506 N_OUT8_Mn8@3506_d N_OUT7_Mn8@3506_g N_VSS_Mn8@3506_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3507 N_OUT8_Mp8@3507_d N_OUT7_Mp8@3507_g N_VDD_Mp8@3507_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3506 N_OUT8_Mp8@3506_d N_OUT7_Mp8@3506_g N_VDD_Mp8@3506_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3505 N_OUT8_Mn8@3505_d N_OUT7_Mn8@3505_g N_VSS_Mn8@3505_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3504 N_OUT8_Mn8@3504_d N_OUT7_Mn8@3504_g N_VSS_Mn8@3504_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3505 N_OUT8_Mp8@3505_d N_OUT7_Mp8@3505_g N_VDD_Mp8@3505_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3504 N_OUT8_Mp8@3504_d N_OUT7_Mp8@3504_g N_VDD_Mp8@3504_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3503 N_OUT8_Mn8@3503_d N_OUT7_Mn8@3503_g N_VSS_Mn8@3503_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3502 N_OUT8_Mn8@3502_d N_OUT7_Mn8@3502_g N_VSS_Mn8@3502_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3503 N_OUT8_Mp8@3503_d N_OUT7_Mp8@3503_g N_VDD_Mp8@3503_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3502 N_OUT8_Mp8@3502_d N_OUT7_Mp8@3502_g N_VDD_Mp8@3502_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3501 N_OUT8_Mn8@3501_d N_OUT7_Mn8@3501_g N_VSS_Mn8@3501_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3500 N_OUT8_Mn8@3500_d N_OUT7_Mn8@3500_g N_VSS_Mn8@3500_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3501 N_OUT8_Mp8@3501_d N_OUT7_Mp8@3501_g N_VDD_Mp8@3501_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3500 N_OUT8_Mp8@3500_d N_OUT7_Mp8@3500_g N_VDD_Mp8@3500_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3499 N_OUT8_Mn8@3499_d N_OUT7_Mn8@3499_g N_VSS_Mn8@3499_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3498 N_OUT8_Mn8@3498_d N_OUT7_Mn8@3498_g N_VSS_Mn8@3498_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3499 N_OUT8_Mp8@3499_d N_OUT7_Mp8@3499_g N_VDD_Mp8@3499_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3498 N_OUT8_Mp8@3498_d N_OUT7_Mp8@3498_g N_VDD_Mp8@3498_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3497 N_OUT8_Mn8@3497_d N_OUT7_Mn8@3497_g N_VSS_Mn8@3497_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3496 N_OUT8_Mn8@3496_d N_OUT7_Mn8@3496_g N_VSS_Mn8@3496_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3497 N_OUT8_Mp8@3497_d N_OUT7_Mp8@3497_g N_VDD_Mp8@3497_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3496 N_OUT8_Mp8@3496_d N_OUT7_Mp8@3496_g N_VDD_Mp8@3496_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3495 N_OUT8_Mn8@3495_d N_OUT7_Mn8@3495_g N_VSS_Mn8@3495_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3494 N_OUT8_Mn8@3494_d N_OUT7_Mn8@3494_g N_VSS_Mn8@3494_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3495 N_OUT8_Mp8@3495_d N_OUT7_Mp8@3495_g N_VDD_Mp8@3495_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3494 N_OUT8_Mp8@3494_d N_OUT7_Mp8@3494_g N_VDD_Mp8@3494_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3493 N_OUT8_Mn8@3493_d N_OUT7_Mn8@3493_g N_VSS_Mn8@3493_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3492 N_OUT8_Mn8@3492_d N_OUT7_Mn8@3492_g N_VSS_Mn8@3492_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3493 N_OUT8_Mp8@3493_d N_OUT7_Mp8@3493_g N_VDD_Mp8@3493_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3492 N_OUT8_Mp8@3492_d N_OUT7_Mp8@3492_g N_VDD_Mp8@3492_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3491 N_OUT8_Mn8@3491_d N_OUT7_Mn8@3491_g N_VSS_Mn8@3491_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3490 N_OUT8_Mn8@3490_d N_OUT7_Mn8@3490_g N_VSS_Mn8@3490_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3491 N_OUT8_Mp8@3491_d N_OUT7_Mp8@3491_g N_VDD_Mp8@3491_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3490 N_OUT8_Mp8@3490_d N_OUT7_Mp8@3490_g N_VDD_Mp8@3490_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3489 N_OUT8_Mn8@3489_d N_OUT7_Mn8@3489_g N_VSS_Mn8@3489_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3488 N_OUT8_Mn8@3488_d N_OUT7_Mn8@3488_g N_VSS_Mn8@3488_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3489 N_OUT8_Mp8@3489_d N_OUT7_Mp8@3489_g N_VDD_Mp8@3489_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3488 N_OUT8_Mp8@3488_d N_OUT7_Mp8@3488_g N_VDD_Mp8@3488_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3487 N_OUT8_Mn8@3487_d N_OUT7_Mn8@3487_g N_VSS_Mn8@3487_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3486 N_OUT8_Mn8@3486_d N_OUT7_Mn8@3486_g N_VSS_Mn8@3486_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3487 N_OUT8_Mp8@3487_d N_OUT7_Mp8@3487_g N_VDD_Mp8@3487_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3486 N_OUT8_Mp8@3486_d N_OUT7_Mp8@3486_g N_VDD_Mp8@3486_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3485 N_OUT8_Mn8@3485_d N_OUT7_Mn8@3485_g N_VSS_Mn8@3485_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3484 N_OUT8_Mn8@3484_d N_OUT7_Mn8@3484_g N_VSS_Mn8@3484_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3485 N_OUT8_Mp8@3485_d N_OUT7_Mp8@3485_g N_VDD_Mp8@3485_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3484 N_OUT8_Mp8@3484_d N_OUT7_Mp8@3484_g N_VDD_Mp8@3484_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3483 N_OUT8_Mn8@3483_d N_OUT7_Mn8@3483_g N_VSS_Mn8@3483_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3482 N_OUT8_Mn8@3482_d N_OUT7_Mn8@3482_g N_VSS_Mn8@3482_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3483 N_OUT8_Mp8@3483_d N_OUT7_Mp8@3483_g N_VDD_Mp8@3483_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3482 N_OUT8_Mp8@3482_d N_OUT7_Mp8@3482_g N_VDD_Mp8@3482_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3481 N_OUT8_Mn8@3481_d N_OUT7_Mn8@3481_g N_VSS_Mn8@3481_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3480 N_OUT8_Mn8@3480_d N_OUT7_Mn8@3480_g N_VSS_Mn8@3480_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3481 N_OUT8_Mp8@3481_d N_OUT7_Mp8@3481_g N_VDD_Mp8@3481_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3480 N_OUT8_Mp8@3480_d N_OUT7_Mp8@3480_g N_VDD_Mp8@3480_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3479 N_OUT8_Mn8@3479_d N_OUT7_Mn8@3479_g N_VSS_Mn8@3479_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3478 N_OUT8_Mn8@3478_d N_OUT7_Mn8@3478_g N_VSS_Mn8@3478_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3479 N_OUT8_Mp8@3479_d N_OUT7_Mp8@3479_g N_VDD_Mp8@3479_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3478 N_OUT8_Mp8@3478_d N_OUT7_Mp8@3478_g N_VDD_Mp8@3478_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3477 N_OUT8_Mn8@3477_d N_OUT7_Mn8@3477_g N_VSS_Mn8@3477_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3476 N_OUT8_Mn8@3476_d N_OUT7_Mn8@3476_g N_VSS_Mn8@3476_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3477 N_OUT8_Mp8@3477_d N_OUT7_Mp8@3477_g N_VDD_Mp8@3477_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3476 N_OUT8_Mp8@3476_d N_OUT7_Mp8@3476_g N_VDD_Mp8@3476_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3475 N_OUT8_Mn8@3475_d N_OUT7_Mn8@3475_g N_VSS_Mn8@3475_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3474 N_OUT8_Mn8@3474_d N_OUT7_Mn8@3474_g N_VSS_Mn8@3474_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3475 N_OUT8_Mp8@3475_d N_OUT7_Mp8@3475_g N_VDD_Mp8@3475_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3474 N_OUT8_Mp8@3474_d N_OUT7_Mp8@3474_g N_VDD_Mp8@3474_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3473 N_OUT8_Mn8@3473_d N_OUT7_Mn8@3473_g N_VSS_Mn8@3473_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3472 N_OUT8_Mn8@3472_d N_OUT7_Mn8@3472_g N_VSS_Mn8@3472_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3473 N_OUT8_Mp8@3473_d N_OUT7_Mp8@3473_g N_VDD_Mp8@3473_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3472 N_OUT8_Mp8@3472_d N_OUT7_Mp8@3472_g N_VDD_Mp8@3472_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3471 N_OUT8_Mn8@3471_d N_OUT7_Mn8@3471_g N_VSS_Mn8@3471_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3470 N_OUT8_Mn8@3470_d N_OUT7_Mn8@3470_g N_VSS_Mn8@3470_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3471 N_OUT8_Mp8@3471_d N_OUT7_Mp8@3471_g N_VDD_Mp8@3471_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3470 N_OUT8_Mp8@3470_d N_OUT7_Mp8@3470_g N_VDD_Mp8@3470_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3469 N_OUT8_Mn8@3469_d N_OUT7_Mn8@3469_g N_VSS_Mn8@3469_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3468 N_OUT8_Mn8@3468_d N_OUT7_Mn8@3468_g N_VSS_Mn8@3468_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3469 N_OUT8_Mp8@3469_d N_OUT7_Mp8@3469_g N_VDD_Mp8@3469_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3468 N_OUT8_Mp8@3468_d N_OUT7_Mp8@3468_g N_VDD_Mp8@3468_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3467 N_OUT8_Mn8@3467_d N_OUT7_Mn8@3467_g N_VSS_Mn8@3467_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3466 N_OUT8_Mn8@3466_d N_OUT7_Mn8@3466_g N_VSS_Mn8@3466_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3467 N_OUT8_Mp8@3467_d N_OUT7_Mp8@3467_g N_VDD_Mp8@3467_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3466 N_OUT8_Mp8@3466_d N_OUT7_Mp8@3466_g N_VDD_Mp8@3466_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3465 N_OUT8_Mn8@3465_d N_OUT7_Mn8@3465_g N_VSS_Mn8@3465_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3464 N_OUT8_Mn8@3464_d N_OUT7_Mn8@3464_g N_VSS_Mn8@3464_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3465 N_OUT8_Mp8@3465_d N_OUT7_Mp8@3465_g N_VDD_Mp8@3465_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3464 N_OUT8_Mp8@3464_d N_OUT7_Mp8@3464_g N_VDD_Mp8@3464_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3463 N_OUT8_Mn8@3463_d N_OUT7_Mn8@3463_g N_VSS_Mn8@3463_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3462 N_OUT8_Mn8@3462_d N_OUT7_Mn8@3462_g N_VSS_Mn8@3462_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3463 N_OUT8_Mp8@3463_d N_OUT7_Mp8@3463_g N_VDD_Mp8@3463_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3462 N_OUT8_Mp8@3462_d N_OUT7_Mp8@3462_g N_VDD_Mp8@3462_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3461 N_OUT8_Mn8@3461_d N_OUT7_Mn8@3461_g N_VSS_Mn8@3461_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3460 N_OUT8_Mn8@3460_d N_OUT7_Mn8@3460_g N_VSS_Mn8@3460_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3461 N_OUT8_Mp8@3461_d N_OUT7_Mp8@3461_g N_VDD_Mp8@3461_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3460 N_OUT8_Mp8@3460_d N_OUT7_Mp8@3460_g N_VDD_Mp8@3460_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3459 N_OUT8_Mn8@3459_d N_OUT7_Mn8@3459_g N_VSS_Mn8@3459_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3458 N_OUT8_Mn8@3458_d N_OUT7_Mn8@3458_g N_VSS_Mn8@3458_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3459 N_OUT8_Mp8@3459_d N_OUT7_Mp8@3459_g N_VDD_Mp8@3459_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3458 N_OUT8_Mp8@3458_d N_OUT7_Mp8@3458_g N_VDD_Mp8@3458_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3457 N_OUT8_Mn8@3457_d N_OUT7_Mn8@3457_g N_VSS_Mn8@3457_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3456 N_OUT8_Mn8@3456_d N_OUT7_Mn8@3456_g N_VSS_Mn8@3456_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3457 N_OUT8_Mp8@3457_d N_OUT7_Mp8@3457_g N_VDD_Mp8@3457_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3456 N_OUT8_Mp8@3456_d N_OUT7_Mp8@3456_g N_VDD_Mp8@3456_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3455 N_OUT8_Mn8@3455_d N_OUT7_Mn8@3455_g N_VSS_Mn8@3455_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3454 N_OUT8_Mn8@3454_d N_OUT7_Mn8@3454_g N_VSS_Mn8@3454_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3455 N_OUT8_Mp8@3455_d N_OUT7_Mp8@3455_g N_VDD_Mp8@3455_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3454 N_OUT8_Mp8@3454_d N_OUT7_Mp8@3454_g N_VDD_Mp8@3454_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3453 N_OUT8_Mn8@3453_d N_OUT7_Mn8@3453_g N_VSS_Mn8@3453_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3452 N_OUT8_Mn8@3452_d N_OUT7_Mn8@3452_g N_VSS_Mn8@3452_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3453 N_OUT8_Mp8@3453_d N_OUT7_Mp8@3453_g N_VDD_Mp8@3453_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3452 N_OUT8_Mp8@3452_d N_OUT7_Mp8@3452_g N_VDD_Mp8@3452_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3451 N_OUT8_Mn8@3451_d N_OUT7_Mn8@3451_g N_VSS_Mn8@3451_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3450 N_OUT8_Mn8@3450_d N_OUT7_Mn8@3450_g N_VSS_Mn8@3450_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3451 N_OUT8_Mp8@3451_d N_OUT7_Mp8@3451_g N_VDD_Mp8@3451_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3450 N_OUT8_Mp8@3450_d N_OUT7_Mp8@3450_g N_VDD_Mp8@3450_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3449 N_OUT8_Mn8@3449_d N_OUT7_Mn8@3449_g N_VSS_Mn8@3449_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3448 N_OUT8_Mn8@3448_d N_OUT7_Mn8@3448_g N_VSS_Mn8@3448_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3449 N_OUT8_Mp8@3449_d N_OUT7_Mp8@3449_g N_VDD_Mp8@3449_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3448 N_OUT8_Mp8@3448_d N_OUT7_Mp8@3448_g N_VDD_Mp8@3448_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3447 N_OUT8_Mn8@3447_d N_OUT7_Mn8@3447_g N_VSS_Mn8@3447_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3446 N_OUT8_Mn8@3446_d N_OUT7_Mn8@3446_g N_VSS_Mn8@3446_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3447 N_OUT8_Mp8@3447_d N_OUT7_Mp8@3447_g N_VDD_Mp8@3447_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3446 N_OUT8_Mp8@3446_d N_OUT7_Mp8@3446_g N_VDD_Mp8@3446_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3445 N_OUT8_Mn8@3445_d N_OUT7_Mn8@3445_g N_VSS_Mn8@3445_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3444 N_OUT8_Mn8@3444_d N_OUT7_Mn8@3444_g N_VSS_Mn8@3444_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3445 N_OUT8_Mp8@3445_d N_OUT7_Mp8@3445_g N_VDD_Mp8@3445_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3444 N_OUT8_Mp8@3444_d N_OUT7_Mp8@3444_g N_VDD_Mp8@3444_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3443 N_OUT8_Mn8@3443_d N_OUT7_Mn8@3443_g N_VSS_Mn8@3443_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3442 N_OUT8_Mn8@3442_d N_OUT7_Mn8@3442_g N_VSS_Mn8@3442_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3443 N_OUT8_Mp8@3443_d N_OUT7_Mp8@3443_g N_VDD_Mp8@3443_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3442 N_OUT8_Mp8@3442_d N_OUT7_Mp8@3442_g N_VDD_Mp8@3442_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3441 N_OUT8_Mn8@3441_d N_OUT7_Mn8@3441_g N_VSS_Mn8@3441_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3440 N_OUT8_Mn8@3440_d N_OUT7_Mn8@3440_g N_VSS_Mn8@3440_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3441 N_OUT8_Mp8@3441_d N_OUT7_Mp8@3441_g N_VDD_Mp8@3441_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3440 N_OUT8_Mp8@3440_d N_OUT7_Mp8@3440_g N_VDD_Mp8@3440_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3439 N_OUT8_Mn8@3439_d N_OUT7_Mn8@3439_g N_VSS_Mn8@3439_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3438 N_OUT8_Mn8@3438_d N_OUT7_Mn8@3438_g N_VSS_Mn8@3438_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3439 N_OUT8_Mp8@3439_d N_OUT7_Mp8@3439_g N_VDD_Mp8@3439_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3438 N_OUT8_Mp8@3438_d N_OUT7_Mp8@3438_g N_VDD_Mp8@3438_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3437 N_OUT8_Mn8@3437_d N_OUT7_Mn8@3437_g N_VSS_Mn8@3437_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3436 N_OUT8_Mn8@3436_d N_OUT7_Mn8@3436_g N_VSS_Mn8@3436_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3437 N_OUT8_Mp8@3437_d N_OUT7_Mp8@3437_g N_VDD_Mp8@3437_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3436 N_OUT8_Mp8@3436_d N_OUT7_Mp8@3436_g N_VDD_Mp8@3436_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3435 N_OUT8_Mn8@3435_d N_OUT7_Mn8@3435_g N_VSS_Mn8@3435_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3434 N_OUT8_Mn8@3434_d N_OUT7_Mn8@3434_g N_VSS_Mn8@3434_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3435 N_OUT8_Mp8@3435_d N_OUT7_Mp8@3435_g N_VDD_Mp8@3435_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3434 N_OUT8_Mp8@3434_d N_OUT7_Mp8@3434_g N_VDD_Mp8@3434_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3433 N_OUT8_Mn8@3433_d N_OUT7_Mn8@3433_g N_VSS_Mn8@3433_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3432 N_OUT8_Mn8@3432_d N_OUT7_Mn8@3432_g N_VSS_Mn8@3432_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3433 N_OUT8_Mp8@3433_d N_OUT7_Mp8@3433_g N_VDD_Mp8@3433_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3432 N_OUT8_Mp8@3432_d N_OUT7_Mp8@3432_g N_VDD_Mp8@3432_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3431 N_OUT8_Mn8@3431_d N_OUT7_Mn8@3431_g N_VSS_Mn8@3431_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3430 N_OUT8_Mn8@3430_d N_OUT7_Mn8@3430_g N_VSS_Mn8@3430_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3431 N_OUT8_Mp8@3431_d N_OUT7_Mp8@3431_g N_VDD_Mp8@3431_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3430 N_OUT8_Mp8@3430_d N_OUT7_Mp8@3430_g N_VDD_Mp8@3430_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3429 N_OUT8_Mn8@3429_d N_OUT7_Mn8@3429_g N_VSS_Mn8@3429_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3428 N_OUT8_Mn8@3428_d N_OUT7_Mn8@3428_g N_VSS_Mn8@3428_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3429 N_OUT8_Mp8@3429_d N_OUT7_Mp8@3429_g N_VDD_Mp8@3429_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3428 N_OUT8_Mp8@3428_d N_OUT7_Mp8@3428_g N_VDD_Mp8@3428_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3427 N_OUT8_Mn8@3427_d N_OUT7_Mn8@3427_g N_VSS_Mn8@3427_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3426 N_OUT8_Mn8@3426_d N_OUT7_Mn8@3426_g N_VSS_Mn8@3426_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3427 N_OUT8_Mp8@3427_d N_OUT7_Mp8@3427_g N_VDD_Mp8@3427_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3426 N_OUT8_Mp8@3426_d N_OUT7_Mp8@3426_g N_VDD_Mp8@3426_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3425 N_OUT8_Mn8@3425_d N_OUT7_Mn8@3425_g N_VSS_Mn8@3425_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3424 N_OUT8_Mn8@3424_d N_OUT7_Mn8@3424_g N_VSS_Mn8@3424_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3425 N_OUT8_Mp8@3425_d N_OUT7_Mp8@3425_g N_VDD_Mp8@3425_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3424 N_OUT8_Mp8@3424_d N_OUT7_Mp8@3424_g N_VDD_Mp8@3424_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3423 N_OUT8_Mn8@3423_d N_OUT7_Mn8@3423_g N_VSS_Mn8@3423_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3422 N_OUT8_Mn8@3422_d N_OUT7_Mn8@3422_g N_VSS_Mn8@3422_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3423 N_OUT8_Mp8@3423_d N_OUT7_Mp8@3423_g N_VDD_Mp8@3423_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3422 N_OUT8_Mp8@3422_d N_OUT7_Mp8@3422_g N_VDD_Mp8@3422_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3421 N_OUT8_Mn8@3421_d N_OUT7_Mn8@3421_g N_VSS_Mn8@3421_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3420 N_OUT8_Mn8@3420_d N_OUT7_Mn8@3420_g N_VSS_Mn8@3420_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3421 N_OUT8_Mp8@3421_d N_OUT7_Mp8@3421_g N_VDD_Mp8@3421_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3420 N_OUT8_Mp8@3420_d N_OUT7_Mp8@3420_g N_VDD_Mp8@3420_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3419 N_OUT8_Mn8@3419_d N_OUT7_Mn8@3419_g N_VSS_Mn8@3419_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3418 N_OUT8_Mn8@3418_d N_OUT7_Mn8@3418_g N_VSS_Mn8@3418_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3419 N_OUT8_Mp8@3419_d N_OUT7_Mp8@3419_g N_VDD_Mp8@3419_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3418 N_OUT8_Mp8@3418_d N_OUT7_Mp8@3418_g N_VDD_Mp8@3418_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3417 N_OUT8_Mn8@3417_d N_OUT7_Mn8@3417_g N_VSS_Mn8@3417_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3416 N_OUT8_Mn8@3416_d N_OUT7_Mn8@3416_g N_VSS_Mn8@3416_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3417 N_OUT8_Mp8@3417_d N_OUT7_Mp8@3417_g N_VDD_Mp8@3417_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3416 N_OUT8_Mp8@3416_d N_OUT7_Mp8@3416_g N_VDD_Mp8@3416_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3415 N_OUT8_Mn8@3415_d N_OUT7_Mn8@3415_g N_VSS_Mn8@3415_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3414 N_OUT8_Mn8@3414_d N_OUT7_Mn8@3414_g N_VSS_Mn8@3414_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3415 N_OUT8_Mp8@3415_d N_OUT7_Mp8@3415_g N_VDD_Mp8@3415_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3414 N_OUT8_Mp8@3414_d N_OUT7_Mp8@3414_g N_VDD_Mp8@3414_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3413 N_OUT8_Mn8@3413_d N_OUT7_Mn8@3413_g N_VSS_Mn8@3413_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3412 N_OUT8_Mn8@3412_d N_OUT7_Mn8@3412_g N_VSS_Mn8@3412_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3413 N_OUT8_Mp8@3413_d N_OUT7_Mp8@3413_g N_VDD_Mp8@3413_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3412 N_OUT8_Mp8@3412_d N_OUT7_Mp8@3412_g N_VDD_Mp8@3412_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3411 N_OUT8_Mn8@3411_d N_OUT7_Mn8@3411_g N_VSS_Mn8@3411_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3410 N_OUT8_Mn8@3410_d N_OUT7_Mn8@3410_g N_VSS_Mn8@3410_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3411 N_OUT8_Mp8@3411_d N_OUT7_Mp8@3411_g N_VDD_Mp8@3411_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3410 N_OUT8_Mp8@3410_d N_OUT7_Mp8@3410_g N_VDD_Mp8@3410_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3409 N_OUT8_Mn8@3409_d N_OUT7_Mn8@3409_g N_VSS_Mn8@3409_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3408 N_OUT8_Mn8@3408_d N_OUT7_Mn8@3408_g N_VSS_Mn8@3408_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3409 N_OUT8_Mp8@3409_d N_OUT7_Mp8@3409_g N_VDD_Mp8@3409_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3408 N_OUT8_Mp8@3408_d N_OUT7_Mp8@3408_g N_VDD_Mp8@3408_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3407 N_OUT8_Mn8@3407_d N_OUT7_Mn8@3407_g N_VSS_Mn8@3407_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3406 N_OUT8_Mn8@3406_d N_OUT7_Mn8@3406_g N_VSS_Mn8@3406_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3407 N_OUT8_Mp8@3407_d N_OUT7_Mp8@3407_g N_VDD_Mp8@3407_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3406 N_OUT8_Mp8@3406_d N_OUT7_Mp8@3406_g N_VDD_Mp8@3406_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3405 N_OUT8_Mn8@3405_d N_OUT7_Mn8@3405_g N_VSS_Mn8@3405_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3404 N_OUT8_Mn8@3404_d N_OUT7_Mn8@3404_g N_VSS_Mn8@3404_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3405 N_OUT8_Mp8@3405_d N_OUT7_Mp8@3405_g N_VDD_Mp8@3405_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3404 N_OUT8_Mp8@3404_d N_OUT7_Mp8@3404_g N_VDD_Mp8@3404_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3403 N_OUT8_Mn8@3403_d N_OUT7_Mn8@3403_g N_VSS_Mn8@3403_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3402 N_OUT8_Mn8@3402_d N_OUT7_Mn8@3402_g N_VSS_Mn8@3402_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3403 N_OUT8_Mp8@3403_d N_OUT7_Mp8@3403_g N_VDD_Mp8@3403_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3402 N_OUT8_Mp8@3402_d N_OUT7_Mp8@3402_g N_VDD_Mp8@3402_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3401 N_OUT8_Mn8@3401_d N_OUT7_Mn8@3401_g N_VSS_Mn8@3401_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3400 N_OUT8_Mn8@3400_d N_OUT7_Mn8@3400_g N_VSS_Mn8@3400_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3401 N_OUT8_Mp8@3401_d N_OUT7_Mp8@3401_g N_VDD_Mp8@3401_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3400 N_OUT8_Mp8@3400_d N_OUT7_Mp8@3400_g N_VDD_Mp8@3400_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3399 N_OUT8_Mn8@3399_d N_OUT7_Mn8@3399_g N_VSS_Mn8@3399_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3398 N_OUT8_Mn8@3398_d N_OUT7_Mn8@3398_g N_VSS_Mn8@3398_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3399 N_OUT8_Mp8@3399_d N_OUT7_Mp8@3399_g N_VDD_Mp8@3399_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3398 N_OUT8_Mp8@3398_d N_OUT7_Mp8@3398_g N_VDD_Mp8@3398_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3397 N_OUT8_Mn8@3397_d N_OUT7_Mn8@3397_g N_VSS_Mn8@3397_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3396 N_OUT8_Mn8@3396_d N_OUT7_Mn8@3396_g N_VSS_Mn8@3396_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3397 N_OUT8_Mp8@3397_d N_OUT7_Mp8@3397_g N_VDD_Mp8@3397_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3396 N_OUT8_Mp8@3396_d N_OUT7_Mp8@3396_g N_VDD_Mp8@3396_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3395 N_OUT8_Mn8@3395_d N_OUT7_Mn8@3395_g N_VSS_Mn8@3395_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3394 N_OUT8_Mn8@3394_d N_OUT7_Mn8@3394_g N_VSS_Mn8@3394_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3395 N_OUT8_Mp8@3395_d N_OUT7_Mp8@3395_g N_VDD_Mp8@3395_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3394 N_OUT8_Mp8@3394_d N_OUT7_Mp8@3394_g N_VDD_Mp8@3394_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3393 N_OUT8_Mn8@3393_d N_OUT7_Mn8@3393_g N_VSS_Mn8@3393_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3392 N_OUT8_Mn8@3392_d N_OUT7_Mn8@3392_g N_VSS_Mn8@3392_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3393 N_OUT8_Mp8@3393_d N_OUT7_Mp8@3393_g N_VDD_Mp8@3393_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3392 N_OUT8_Mp8@3392_d N_OUT7_Mp8@3392_g N_VDD_Mp8@3392_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3391 N_OUT8_Mn8@3391_d N_OUT7_Mn8@3391_g N_VSS_Mn8@3391_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3390 N_OUT8_Mn8@3390_d N_OUT7_Mn8@3390_g N_VSS_Mn8@3390_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3391 N_OUT8_Mp8@3391_d N_OUT7_Mp8@3391_g N_VDD_Mp8@3391_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3390 N_OUT8_Mp8@3390_d N_OUT7_Mp8@3390_g N_VDD_Mp8@3390_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3389 N_OUT8_Mn8@3389_d N_OUT7_Mn8@3389_g N_VSS_Mn8@3389_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3388 N_OUT8_Mn8@3388_d N_OUT7_Mn8@3388_g N_VSS_Mn8@3388_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3389 N_OUT8_Mp8@3389_d N_OUT7_Mp8@3389_g N_VDD_Mp8@3389_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3388 N_OUT8_Mp8@3388_d N_OUT7_Mp8@3388_g N_VDD_Mp8@3388_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3387 N_OUT8_Mn8@3387_d N_OUT7_Mn8@3387_g N_VSS_Mn8@3387_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3386 N_OUT8_Mn8@3386_d N_OUT7_Mn8@3386_g N_VSS_Mn8@3386_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3387 N_OUT8_Mp8@3387_d N_OUT7_Mp8@3387_g N_VDD_Mp8@3387_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3386 N_OUT8_Mp8@3386_d N_OUT7_Mp8@3386_g N_VDD_Mp8@3386_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3385 N_OUT8_Mn8@3385_d N_OUT7_Mn8@3385_g N_VSS_Mn8@3385_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3384 N_OUT8_Mn8@3384_d N_OUT7_Mn8@3384_g N_VSS_Mn8@3384_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3385 N_OUT8_Mp8@3385_d N_OUT7_Mp8@3385_g N_VDD_Mp8@3385_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3384 N_OUT8_Mp8@3384_d N_OUT7_Mp8@3384_g N_VDD_Mp8@3384_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3383 N_OUT8_Mn8@3383_d N_OUT7_Mn8@3383_g N_VSS_Mn8@3383_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3382 N_OUT8_Mn8@3382_d N_OUT7_Mn8@3382_g N_VSS_Mn8@3382_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3383 N_OUT8_Mp8@3383_d N_OUT7_Mp8@3383_g N_VDD_Mp8@3383_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3382 N_OUT8_Mp8@3382_d N_OUT7_Mp8@3382_g N_VDD_Mp8@3382_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3381 N_OUT8_Mn8@3381_d N_OUT7_Mn8@3381_g N_VSS_Mn8@3381_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3380 N_OUT8_Mn8@3380_d N_OUT7_Mn8@3380_g N_VSS_Mn8@3380_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3381 N_OUT8_Mp8@3381_d N_OUT7_Mp8@3381_g N_VDD_Mp8@3381_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3380 N_OUT8_Mp8@3380_d N_OUT7_Mp8@3380_g N_VDD_Mp8@3380_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3379 N_OUT8_Mn8@3379_d N_OUT7_Mn8@3379_g N_VSS_Mn8@3379_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3378 N_OUT8_Mn8@3378_d N_OUT7_Mn8@3378_g N_VSS_Mn8@3378_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3379 N_OUT8_Mp8@3379_d N_OUT7_Mp8@3379_g N_VDD_Mp8@3379_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3378 N_OUT8_Mp8@3378_d N_OUT7_Mp8@3378_g N_VDD_Mp8@3378_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3377 N_OUT8_Mn8@3377_d N_OUT7_Mn8@3377_g N_VSS_Mn8@3377_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3376 N_OUT8_Mn8@3376_d N_OUT7_Mn8@3376_g N_VSS_Mn8@3376_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3377 N_OUT8_Mp8@3377_d N_OUT7_Mp8@3377_g N_VDD_Mp8@3377_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3376 N_OUT8_Mp8@3376_d N_OUT7_Mp8@3376_g N_VDD_Mp8@3376_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3375 N_OUT8_Mn8@3375_d N_OUT7_Mn8@3375_g N_VSS_Mn8@3375_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3374 N_OUT8_Mn8@3374_d N_OUT7_Mn8@3374_g N_VSS_Mn8@3374_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3375 N_OUT8_Mp8@3375_d N_OUT7_Mp8@3375_g N_VDD_Mp8@3375_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3374 N_OUT8_Mp8@3374_d N_OUT7_Mp8@3374_g N_VDD_Mp8@3374_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3373 N_OUT8_Mn8@3373_d N_OUT7_Mn8@3373_g N_VSS_Mn8@3373_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3372 N_OUT8_Mn8@3372_d N_OUT7_Mn8@3372_g N_VSS_Mn8@3372_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3373 N_OUT8_Mp8@3373_d N_OUT7_Mp8@3373_g N_VDD_Mp8@3373_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3372 N_OUT8_Mp8@3372_d N_OUT7_Mp8@3372_g N_VDD_Mp8@3372_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3371 N_OUT8_Mn8@3371_d N_OUT7_Mn8@3371_g N_VSS_Mn8@3371_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3370 N_OUT8_Mn8@3370_d N_OUT7_Mn8@3370_g N_VSS_Mn8@3370_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3371 N_OUT8_Mp8@3371_d N_OUT7_Mp8@3371_g N_VDD_Mp8@3371_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3370 N_OUT8_Mp8@3370_d N_OUT7_Mp8@3370_g N_VDD_Mp8@3370_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3369 N_OUT8_Mn8@3369_d N_OUT7_Mn8@3369_g N_VSS_Mn8@3369_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3368 N_OUT8_Mn8@3368_d N_OUT7_Mn8@3368_g N_VSS_Mn8@3368_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3369 N_OUT8_Mp8@3369_d N_OUT7_Mp8@3369_g N_VDD_Mp8@3369_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3368 N_OUT8_Mp8@3368_d N_OUT7_Mp8@3368_g N_VDD_Mp8@3368_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3367 N_OUT8_Mn8@3367_d N_OUT7_Mn8@3367_g N_VSS_Mn8@3367_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3366 N_OUT8_Mn8@3366_d N_OUT7_Mn8@3366_g N_VSS_Mn8@3366_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3367 N_OUT8_Mp8@3367_d N_OUT7_Mp8@3367_g N_VDD_Mp8@3367_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3366 N_OUT8_Mp8@3366_d N_OUT7_Mp8@3366_g N_VDD_Mp8@3366_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3365 N_OUT8_Mn8@3365_d N_OUT7_Mn8@3365_g N_VSS_Mn8@3365_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3364 N_OUT8_Mn8@3364_d N_OUT7_Mn8@3364_g N_VSS_Mn8@3364_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3365 N_OUT8_Mp8@3365_d N_OUT7_Mp8@3365_g N_VDD_Mp8@3365_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3364 N_OUT8_Mp8@3364_d N_OUT7_Mp8@3364_g N_VDD_Mp8@3364_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3363 N_OUT8_Mn8@3363_d N_OUT7_Mn8@3363_g N_VSS_Mn8@3363_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3362 N_OUT8_Mn8@3362_d N_OUT7_Mn8@3362_g N_VSS_Mn8@3362_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3363 N_OUT8_Mp8@3363_d N_OUT7_Mp8@3363_g N_VDD_Mp8@3363_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3362 N_OUT8_Mp8@3362_d N_OUT7_Mp8@3362_g N_VDD_Mp8@3362_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3361 N_OUT8_Mn8@3361_d N_OUT7_Mn8@3361_g N_VSS_Mn8@3361_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3360 N_OUT8_Mn8@3360_d N_OUT7_Mn8@3360_g N_VSS_Mn8@3360_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3361 N_OUT8_Mp8@3361_d N_OUT7_Mp8@3361_g N_VDD_Mp8@3361_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3360 N_OUT8_Mp8@3360_d N_OUT7_Mp8@3360_g N_VDD_Mp8@3360_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3359 N_OUT8_Mn8@3359_d N_OUT7_Mn8@3359_g N_VSS_Mn8@3359_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3358 N_OUT8_Mn8@3358_d N_OUT7_Mn8@3358_g N_VSS_Mn8@3358_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3359 N_OUT8_Mp8@3359_d N_OUT7_Mp8@3359_g N_VDD_Mp8@3359_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3358 N_OUT8_Mp8@3358_d N_OUT7_Mp8@3358_g N_VDD_Mp8@3358_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3357 N_OUT8_Mn8@3357_d N_OUT7_Mn8@3357_g N_VSS_Mn8@3357_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3356 N_OUT8_Mn8@3356_d N_OUT7_Mn8@3356_g N_VSS_Mn8@3356_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3357 N_OUT8_Mp8@3357_d N_OUT7_Mp8@3357_g N_VDD_Mp8@3357_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3356 N_OUT8_Mp8@3356_d N_OUT7_Mp8@3356_g N_VDD_Mp8@3356_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3355 N_OUT8_Mn8@3355_d N_OUT7_Mn8@3355_g N_VSS_Mn8@3355_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3354 N_OUT8_Mn8@3354_d N_OUT7_Mn8@3354_g N_VSS_Mn8@3354_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3355 N_OUT8_Mp8@3355_d N_OUT7_Mp8@3355_g N_VDD_Mp8@3355_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3354 N_OUT8_Mp8@3354_d N_OUT7_Mp8@3354_g N_VDD_Mp8@3354_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3353 N_OUT8_Mn8@3353_d N_OUT7_Mn8@3353_g N_VSS_Mn8@3353_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3352 N_OUT8_Mn8@3352_d N_OUT7_Mn8@3352_g N_VSS_Mn8@3352_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3353 N_OUT8_Mp8@3353_d N_OUT7_Mp8@3353_g N_VDD_Mp8@3353_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3352 N_OUT8_Mp8@3352_d N_OUT7_Mp8@3352_g N_VDD_Mp8@3352_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3351 N_OUT8_Mn8@3351_d N_OUT7_Mn8@3351_g N_VSS_Mn8@3351_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3350 N_OUT8_Mn8@3350_d N_OUT7_Mn8@3350_g N_VSS_Mn8@3350_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3351 N_OUT8_Mp8@3351_d N_OUT7_Mp8@3351_g N_VDD_Mp8@3351_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3350 N_OUT8_Mp8@3350_d N_OUT7_Mp8@3350_g N_VDD_Mp8@3350_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3349 N_OUT8_Mn8@3349_d N_OUT7_Mn8@3349_g N_VSS_Mn8@3349_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3348 N_OUT8_Mn8@3348_d N_OUT7_Mn8@3348_g N_VSS_Mn8@3348_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3349 N_OUT8_Mp8@3349_d N_OUT7_Mp8@3349_g N_VDD_Mp8@3349_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3348 N_OUT8_Mp8@3348_d N_OUT7_Mp8@3348_g N_VDD_Mp8@3348_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3347 N_OUT8_Mn8@3347_d N_OUT7_Mn8@3347_g N_VSS_Mn8@3347_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3346 N_OUT8_Mn8@3346_d N_OUT7_Mn8@3346_g N_VSS_Mn8@3346_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3347 N_OUT8_Mp8@3347_d N_OUT7_Mp8@3347_g N_VDD_Mp8@3347_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3346 N_OUT8_Mp8@3346_d N_OUT7_Mp8@3346_g N_VDD_Mp8@3346_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3345 N_OUT8_Mn8@3345_d N_OUT7_Mn8@3345_g N_VSS_Mn8@3345_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3344 N_OUT8_Mn8@3344_d N_OUT7_Mn8@3344_g N_VSS_Mn8@3344_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3345 N_OUT8_Mp8@3345_d N_OUT7_Mp8@3345_g N_VDD_Mp8@3345_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3344 N_OUT8_Mp8@3344_d N_OUT7_Mp8@3344_g N_VDD_Mp8@3344_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3343 N_OUT8_Mn8@3343_d N_OUT7_Mn8@3343_g N_VSS_Mn8@3343_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3342 N_OUT8_Mn8@3342_d N_OUT7_Mn8@3342_g N_VSS_Mn8@3342_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3343 N_OUT8_Mp8@3343_d N_OUT7_Mp8@3343_g N_VDD_Mp8@3343_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3342 N_OUT8_Mp8@3342_d N_OUT7_Mp8@3342_g N_VDD_Mp8@3342_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3341 N_OUT8_Mn8@3341_d N_OUT7_Mn8@3341_g N_VSS_Mn8@3341_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3340 N_OUT8_Mn8@3340_d N_OUT7_Mn8@3340_g N_VSS_Mn8@3340_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3341 N_OUT8_Mp8@3341_d N_OUT7_Mp8@3341_g N_VDD_Mp8@3341_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3340 N_OUT8_Mp8@3340_d N_OUT7_Mp8@3340_g N_VDD_Mp8@3340_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3339 N_OUT8_Mn8@3339_d N_OUT7_Mn8@3339_g N_VSS_Mn8@3339_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3338 N_OUT8_Mn8@3338_d N_OUT7_Mn8@3338_g N_VSS_Mn8@3338_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3339 N_OUT8_Mp8@3339_d N_OUT7_Mp8@3339_g N_VDD_Mp8@3339_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3338 N_OUT8_Mp8@3338_d N_OUT7_Mp8@3338_g N_VDD_Mp8@3338_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3337 N_OUT8_Mn8@3337_d N_OUT7_Mn8@3337_g N_VSS_Mn8@3337_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3336 N_OUT8_Mn8@3336_d N_OUT7_Mn8@3336_g N_VSS_Mn8@3336_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3337 N_OUT8_Mp8@3337_d N_OUT7_Mp8@3337_g N_VDD_Mp8@3337_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3336 N_OUT8_Mp8@3336_d N_OUT7_Mp8@3336_g N_VDD_Mp8@3336_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3335 N_OUT8_Mn8@3335_d N_OUT7_Mn8@3335_g N_VSS_Mn8@3335_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3334 N_OUT8_Mn8@3334_d N_OUT7_Mn8@3334_g N_VSS_Mn8@3334_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3335 N_OUT8_Mp8@3335_d N_OUT7_Mp8@3335_g N_VDD_Mp8@3335_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3334 N_OUT8_Mp8@3334_d N_OUT7_Mp8@3334_g N_VDD_Mp8@3334_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3333 N_OUT8_Mn8@3333_d N_OUT7_Mn8@3333_g N_VSS_Mn8@3333_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3332 N_OUT8_Mn8@3332_d N_OUT7_Mn8@3332_g N_VSS_Mn8@3332_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3333 N_OUT8_Mp8@3333_d N_OUT7_Mp8@3333_g N_VDD_Mp8@3333_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3332 N_OUT8_Mp8@3332_d N_OUT7_Mp8@3332_g N_VDD_Mp8@3332_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3331 N_OUT8_Mn8@3331_d N_OUT7_Mn8@3331_g N_VSS_Mn8@3331_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3330 N_OUT8_Mn8@3330_d N_OUT7_Mn8@3330_g N_VSS_Mn8@3330_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3331 N_OUT8_Mp8@3331_d N_OUT7_Mp8@3331_g N_VDD_Mp8@3331_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3330 N_OUT8_Mp8@3330_d N_OUT7_Mp8@3330_g N_VDD_Mp8@3330_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3329 N_OUT8_Mn8@3329_d N_OUT7_Mn8@3329_g N_VSS_Mn8@3329_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3328 N_OUT8_Mn8@3328_d N_OUT7_Mn8@3328_g N_VSS_Mn8@3328_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3329 N_OUT8_Mp8@3329_d N_OUT7_Mp8@3329_g N_VDD_Mp8@3329_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3328 N_OUT8_Mp8@3328_d N_OUT7_Mp8@3328_g N_VDD_Mp8@3328_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3327 N_OUT8_Mn8@3327_d N_OUT7_Mn8@3327_g N_VSS_Mn8@3327_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3326 N_OUT8_Mn8@3326_d N_OUT7_Mn8@3326_g N_VSS_Mn8@3326_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3327 N_OUT8_Mp8@3327_d N_OUT7_Mp8@3327_g N_VDD_Mp8@3327_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3326 N_OUT8_Mp8@3326_d N_OUT7_Mp8@3326_g N_VDD_Mp8@3326_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3325 N_OUT8_Mn8@3325_d N_OUT7_Mn8@3325_g N_VSS_Mn8@3325_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3324 N_OUT8_Mn8@3324_d N_OUT7_Mn8@3324_g N_VSS_Mn8@3324_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3325 N_OUT8_Mp8@3325_d N_OUT7_Mp8@3325_g N_VDD_Mp8@3325_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3324 N_OUT8_Mp8@3324_d N_OUT7_Mp8@3324_g N_VDD_Mp8@3324_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3323 N_OUT8_Mn8@3323_d N_OUT7_Mn8@3323_g N_VSS_Mn8@3323_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3322 N_OUT8_Mn8@3322_d N_OUT7_Mn8@3322_g N_VSS_Mn8@3322_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3323 N_OUT8_Mp8@3323_d N_OUT7_Mp8@3323_g N_VDD_Mp8@3323_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3322 N_OUT8_Mp8@3322_d N_OUT7_Mp8@3322_g N_VDD_Mp8@3322_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3321 N_OUT8_Mn8@3321_d N_OUT7_Mn8@3321_g N_VSS_Mn8@3321_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3320 N_OUT8_Mn8@3320_d N_OUT7_Mn8@3320_g N_VSS_Mn8@3320_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3321 N_OUT8_Mp8@3321_d N_OUT7_Mp8@3321_g N_VDD_Mp8@3321_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3320 N_OUT8_Mp8@3320_d N_OUT7_Mp8@3320_g N_VDD_Mp8@3320_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3319 N_OUT8_Mn8@3319_d N_OUT7_Mn8@3319_g N_VSS_Mn8@3319_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3318 N_OUT8_Mn8@3318_d N_OUT7_Mn8@3318_g N_VSS_Mn8@3318_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3319 N_OUT8_Mp8@3319_d N_OUT7_Mp8@3319_g N_VDD_Mp8@3319_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3318 N_OUT8_Mp8@3318_d N_OUT7_Mp8@3318_g N_VDD_Mp8@3318_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3317 N_OUT8_Mn8@3317_d N_OUT7_Mn8@3317_g N_VSS_Mn8@3317_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3316 N_OUT8_Mn8@3316_d N_OUT7_Mn8@3316_g N_VSS_Mn8@3316_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3317 N_OUT8_Mp8@3317_d N_OUT7_Mp8@3317_g N_VDD_Mp8@3317_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3316 N_OUT8_Mp8@3316_d N_OUT7_Mp8@3316_g N_VDD_Mp8@3316_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3315 N_OUT8_Mn8@3315_d N_OUT7_Mn8@3315_g N_VSS_Mn8@3315_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3314 N_OUT8_Mn8@3314_d N_OUT7_Mn8@3314_g N_VSS_Mn8@3314_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3315 N_OUT8_Mp8@3315_d N_OUT7_Mp8@3315_g N_VDD_Mp8@3315_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3314 N_OUT8_Mp8@3314_d N_OUT7_Mp8@3314_g N_VDD_Mp8@3314_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3313 N_OUT8_Mn8@3313_d N_OUT7_Mn8@3313_g N_VSS_Mn8@3313_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3312 N_OUT8_Mn8@3312_d N_OUT7_Mn8@3312_g N_VSS_Mn8@3312_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3313 N_OUT8_Mp8@3313_d N_OUT7_Mp8@3313_g N_VDD_Mp8@3313_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3312 N_OUT8_Mp8@3312_d N_OUT7_Mp8@3312_g N_VDD_Mp8@3312_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3311 N_OUT8_Mn8@3311_d N_OUT7_Mn8@3311_g N_VSS_Mn8@3311_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3310 N_OUT8_Mn8@3310_d N_OUT7_Mn8@3310_g N_VSS_Mn8@3310_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3311 N_OUT8_Mp8@3311_d N_OUT7_Mp8@3311_g N_VDD_Mp8@3311_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3310 N_OUT8_Mp8@3310_d N_OUT7_Mp8@3310_g N_VDD_Mp8@3310_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3309 N_OUT8_Mn8@3309_d N_OUT7_Mn8@3309_g N_VSS_Mn8@3309_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3308 N_OUT8_Mn8@3308_d N_OUT7_Mn8@3308_g N_VSS_Mn8@3308_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3309 N_OUT8_Mp8@3309_d N_OUT7_Mp8@3309_g N_VDD_Mp8@3309_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3308 N_OUT8_Mp8@3308_d N_OUT7_Mp8@3308_g N_VDD_Mp8@3308_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3307 N_OUT8_Mn8@3307_d N_OUT7_Mn8@3307_g N_VSS_Mn8@3307_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3306 N_OUT8_Mn8@3306_d N_OUT7_Mn8@3306_g N_VSS_Mn8@3306_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3307 N_OUT8_Mp8@3307_d N_OUT7_Mp8@3307_g N_VDD_Mp8@3307_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3306 N_OUT8_Mp8@3306_d N_OUT7_Mp8@3306_g N_VDD_Mp8@3306_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3305 N_OUT8_Mn8@3305_d N_OUT7_Mn8@3305_g N_VSS_Mn8@3305_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3304 N_OUT8_Mn8@3304_d N_OUT7_Mn8@3304_g N_VSS_Mn8@3304_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3305 N_OUT8_Mp8@3305_d N_OUT7_Mp8@3305_g N_VDD_Mp8@3305_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3304 N_OUT8_Mp8@3304_d N_OUT7_Mp8@3304_g N_VDD_Mp8@3304_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3303 N_OUT8_Mn8@3303_d N_OUT7_Mn8@3303_g N_VSS_Mn8@3303_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3302 N_OUT8_Mn8@3302_d N_OUT7_Mn8@3302_g N_VSS_Mn8@3302_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3303 N_OUT8_Mp8@3303_d N_OUT7_Mp8@3303_g N_VDD_Mp8@3303_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3302 N_OUT8_Mp8@3302_d N_OUT7_Mp8@3302_g N_VDD_Mp8@3302_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3301 N_OUT8_Mn8@3301_d N_OUT7_Mn8@3301_g N_VSS_Mn8@3301_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3300 N_OUT8_Mn8@3300_d N_OUT7_Mn8@3300_g N_VSS_Mn8@3300_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3301 N_OUT8_Mp8@3301_d N_OUT7_Mp8@3301_g N_VDD_Mp8@3301_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3300 N_OUT8_Mp8@3300_d N_OUT7_Mp8@3300_g N_VDD_Mp8@3300_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3299 N_OUT8_Mn8@3299_d N_OUT7_Mn8@3299_g N_VSS_Mn8@3299_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3298 N_OUT8_Mn8@3298_d N_OUT7_Mn8@3298_g N_VSS_Mn8@3298_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3299 N_OUT8_Mp8@3299_d N_OUT7_Mp8@3299_g N_VDD_Mp8@3299_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3298 N_OUT8_Mp8@3298_d N_OUT7_Mp8@3298_g N_VDD_Mp8@3298_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3297 N_OUT8_Mn8@3297_d N_OUT7_Mn8@3297_g N_VSS_Mn8@3297_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3296 N_OUT8_Mn8@3296_d N_OUT7_Mn8@3296_g N_VSS_Mn8@3296_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3297 N_OUT8_Mp8@3297_d N_OUT7_Mp8@3297_g N_VDD_Mp8@3297_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3296 N_OUT8_Mp8@3296_d N_OUT7_Mp8@3296_g N_VDD_Mp8@3296_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3295 N_OUT8_Mn8@3295_d N_OUT7_Mn8@3295_g N_VSS_Mn8@3295_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3294 N_OUT8_Mn8@3294_d N_OUT7_Mn8@3294_g N_VSS_Mn8@3294_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3295 N_OUT8_Mp8@3295_d N_OUT7_Mp8@3295_g N_VDD_Mp8@3295_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3294 N_OUT8_Mp8@3294_d N_OUT7_Mp8@3294_g N_VDD_Mp8@3294_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3293 N_OUT8_Mn8@3293_d N_OUT7_Mn8@3293_g N_VSS_Mn8@3293_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3292 N_OUT8_Mn8@3292_d N_OUT7_Mn8@3292_g N_VSS_Mn8@3292_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3293 N_OUT8_Mp8@3293_d N_OUT7_Mp8@3293_g N_VDD_Mp8@3293_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3292 N_OUT8_Mp8@3292_d N_OUT7_Mp8@3292_g N_VDD_Mp8@3292_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3291 N_OUT8_Mn8@3291_d N_OUT7_Mn8@3291_g N_VSS_Mn8@3291_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3290 N_OUT8_Mn8@3290_d N_OUT7_Mn8@3290_g N_VSS_Mn8@3290_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3291 N_OUT8_Mp8@3291_d N_OUT7_Mp8@3291_g N_VDD_Mp8@3291_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3290 N_OUT8_Mp8@3290_d N_OUT7_Mp8@3290_g N_VDD_Mp8@3290_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3289 N_OUT8_Mn8@3289_d N_OUT7_Mn8@3289_g N_VSS_Mn8@3289_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3288 N_OUT8_Mn8@3288_d N_OUT7_Mn8@3288_g N_VSS_Mn8@3288_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3289 N_OUT8_Mp8@3289_d N_OUT7_Mp8@3289_g N_VDD_Mp8@3289_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3288 N_OUT8_Mp8@3288_d N_OUT7_Mp8@3288_g N_VDD_Mp8@3288_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3287 N_OUT8_Mn8@3287_d N_OUT7_Mn8@3287_g N_VSS_Mn8@3287_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3286 N_OUT8_Mn8@3286_d N_OUT7_Mn8@3286_g N_VSS_Mn8@3286_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3287 N_OUT8_Mp8@3287_d N_OUT7_Mp8@3287_g N_VDD_Mp8@3287_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3286 N_OUT8_Mp8@3286_d N_OUT7_Mp8@3286_g N_VDD_Mp8@3286_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3285 N_OUT8_Mn8@3285_d N_OUT7_Mn8@3285_g N_VSS_Mn8@3285_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3284 N_OUT8_Mn8@3284_d N_OUT7_Mn8@3284_g N_VSS_Mn8@3284_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3285 N_OUT8_Mp8@3285_d N_OUT7_Mp8@3285_g N_VDD_Mp8@3285_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3284 N_OUT8_Mp8@3284_d N_OUT7_Mp8@3284_g N_VDD_Mp8@3284_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3283 N_OUT8_Mn8@3283_d N_OUT7_Mn8@3283_g N_VSS_Mn8@3283_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3282 N_OUT8_Mn8@3282_d N_OUT7_Mn8@3282_g N_VSS_Mn8@3282_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3283 N_OUT8_Mp8@3283_d N_OUT7_Mp8@3283_g N_VDD_Mp8@3283_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3282 N_OUT8_Mp8@3282_d N_OUT7_Mp8@3282_g N_VDD_Mp8@3282_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3281 N_OUT8_Mn8@3281_d N_OUT7_Mn8@3281_g N_VSS_Mn8@3281_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3280 N_OUT8_Mn8@3280_d N_OUT7_Mn8@3280_g N_VSS_Mn8@3280_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3281 N_OUT8_Mp8@3281_d N_OUT7_Mp8@3281_g N_VDD_Mp8@3281_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3280 N_OUT8_Mp8@3280_d N_OUT7_Mp8@3280_g N_VDD_Mp8@3280_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3279 N_OUT8_Mn8@3279_d N_OUT7_Mn8@3279_g N_VSS_Mn8@3279_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3278 N_OUT8_Mn8@3278_d N_OUT7_Mn8@3278_g N_VSS_Mn8@3278_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3279 N_OUT8_Mp8@3279_d N_OUT7_Mp8@3279_g N_VDD_Mp8@3279_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3278 N_OUT8_Mp8@3278_d N_OUT7_Mp8@3278_g N_VDD_Mp8@3278_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3277 N_OUT8_Mn8@3277_d N_OUT7_Mn8@3277_g N_VSS_Mn8@3277_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3276 N_OUT8_Mn8@3276_d N_OUT7_Mn8@3276_g N_VSS_Mn8@3276_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3277 N_OUT8_Mp8@3277_d N_OUT7_Mp8@3277_g N_VDD_Mp8@3277_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3276 N_OUT8_Mp8@3276_d N_OUT7_Mp8@3276_g N_VDD_Mp8@3276_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3275 N_OUT8_Mn8@3275_d N_OUT7_Mn8@3275_g N_VSS_Mn8@3275_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3274 N_OUT8_Mn8@3274_d N_OUT7_Mn8@3274_g N_VSS_Mn8@3274_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3275 N_OUT8_Mp8@3275_d N_OUT7_Mp8@3275_g N_VDD_Mp8@3275_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3274 N_OUT8_Mp8@3274_d N_OUT7_Mp8@3274_g N_VDD_Mp8@3274_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3273 N_OUT8_Mn8@3273_d N_OUT7_Mn8@3273_g N_VSS_Mn8@3273_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3272 N_OUT8_Mn8@3272_d N_OUT7_Mn8@3272_g N_VSS_Mn8@3272_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3273 N_OUT8_Mp8@3273_d N_OUT7_Mp8@3273_g N_VDD_Mp8@3273_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3272 N_OUT8_Mp8@3272_d N_OUT7_Mp8@3272_g N_VDD_Mp8@3272_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3271 N_OUT8_Mn8@3271_d N_OUT7_Mn8@3271_g N_VSS_Mn8@3271_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3270 N_OUT8_Mn8@3270_d N_OUT7_Mn8@3270_g N_VSS_Mn8@3270_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3271 N_OUT8_Mp8@3271_d N_OUT7_Mp8@3271_g N_VDD_Mp8@3271_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3270 N_OUT8_Mp8@3270_d N_OUT7_Mp8@3270_g N_VDD_Mp8@3270_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3269 N_OUT8_Mn8@3269_d N_OUT7_Mn8@3269_g N_VSS_Mn8@3269_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3268 N_OUT8_Mn8@3268_d N_OUT7_Mn8@3268_g N_VSS_Mn8@3268_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3269 N_OUT8_Mp8@3269_d N_OUT7_Mp8@3269_g N_VDD_Mp8@3269_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3268 N_OUT8_Mp8@3268_d N_OUT7_Mp8@3268_g N_VDD_Mp8@3268_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3267 N_OUT8_Mn8@3267_d N_OUT7_Mn8@3267_g N_VSS_Mn8@3267_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3266 N_OUT8_Mn8@3266_d N_OUT7_Mn8@3266_g N_VSS_Mn8@3266_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3267 N_OUT8_Mp8@3267_d N_OUT7_Mp8@3267_g N_VDD_Mp8@3267_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3266 N_OUT8_Mp8@3266_d N_OUT7_Mp8@3266_g N_VDD_Mp8@3266_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3265 N_OUT8_Mn8@3265_d N_OUT7_Mn8@3265_g N_VSS_Mn8@3265_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3264 N_OUT8_Mn8@3264_d N_OUT7_Mn8@3264_g N_VSS_Mn8@3264_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3265 N_OUT8_Mp8@3265_d N_OUT7_Mp8@3265_g N_VDD_Mp8@3265_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3264 N_OUT8_Mp8@3264_d N_OUT7_Mp8@3264_g N_VDD_Mp8@3264_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3263 N_OUT8_Mn8@3263_d N_OUT7_Mn8@3263_g N_VSS_Mn8@3263_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3262 N_OUT8_Mn8@3262_d N_OUT7_Mn8@3262_g N_VSS_Mn8@3262_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3263 N_OUT8_Mp8@3263_d N_OUT7_Mp8@3263_g N_VDD_Mp8@3263_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3262 N_OUT8_Mp8@3262_d N_OUT7_Mp8@3262_g N_VDD_Mp8@3262_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3261 N_OUT8_Mn8@3261_d N_OUT7_Mn8@3261_g N_VSS_Mn8@3261_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3260 N_OUT8_Mn8@3260_d N_OUT7_Mn8@3260_g N_VSS_Mn8@3260_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3261 N_OUT8_Mp8@3261_d N_OUT7_Mp8@3261_g N_VDD_Mp8@3261_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3260 N_OUT8_Mp8@3260_d N_OUT7_Mp8@3260_g N_VDD_Mp8@3260_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3259 N_OUT8_Mn8@3259_d N_OUT7_Mn8@3259_g N_VSS_Mn8@3259_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3258 N_OUT8_Mn8@3258_d N_OUT7_Mn8@3258_g N_VSS_Mn8@3258_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3259 N_OUT8_Mp8@3259_d N_OUT7_Mp8@3259_g N_VDD_Mp8@3259_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3258 N_OUT8_Mp8@3258_d N_OUT7_Mp8@3258_g N_VDD_Mp8@3258_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3257 N_OUT8_Mn8@3257_d N_OUT7_Mn8@3257_g N_VSS_Mn8@3257_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3256 N_OUT8_Mn8@3256_d N_OUT7_Mn8@3256_g N_VSS_Mn8@3256_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3257 N_OUT8_Mp8@3257_d N_OUT7_Mp8@3257_g N_VDD_Mp8@3257_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3256 N_OUT8_Mp8@3256_d N_OUT7_Mp8@3256_g N_VDD_Mp8@3256_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3255 N_OUT8_Mn8@3255_d N_OUT7_Mn8@3255_g N_VSS_Mn8@3255_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3254 N_OUT8_Mn8@3254_d N_OUT7_Mn8@3254_g N_VSS_Mn8@3254_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3255 N_OUT8_Mp8@3255_d N_OUT7_Mp8@3255_g N_VDD_Mp8@3255_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3254 N_OUT8_Mp8@3254_d N_OUT7_Mp8@3254_g N_VDD_Mp8@3254_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3253 N_OUT8_Mn8@3253_d N_OUT7_Mn8@3253_g N_VSS_Mn8@3253_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3252 N_OUT8_Mn8@3252_d N_OUT7_Mn8@3252_g N_VSS_Mn8@3252_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3253 N_OUT8_Mp8@3253_d N_OUT7_Mp8@3253_g N_VDD_Mp8@3253_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3252 N_OUT8_Mp8@3252_d N_OUT7_Mp8@3252_g N_VDD_Mp8@3252_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3251 N_OUT8_Mn8@3251_d N_OUT7_Mn8@3251_g N_VSS_Mn8@3251_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3250 N_OUT8_Mn8@3250_d N_OUT7_Mn8@3250_g N_VSS_Mn8@3250_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3251 N_OUT8_Mp8@3251_d N_OUT7_Mp8@3251_g N_VDD_Mp8@3251_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3250 N_OUT8_Mp8@3250_d N_OUT7_Mp8@3250_g N_VDD_Mp8@3250_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3249 N_OUT8_Mn8@3249_d N_OUT7_Mn8@3249_g N_VSS_Mn8@3249_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3248 N_OUT8_Mn8@3248_d N_OUT7_Mn8@3248_g N_VSS_Mn8@3248_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3249 N_OUT8_Mp8@3249_d N_OUT7_Mp8@3249_g N_VDD_Mp8@3249_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3248 N_OUT8_Mp8@3248_d N_OUT7_Mp8@3248_g N_VDD_Mp8@3248_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3247 N_OUT8_Mn8@3247_d N_OUT7_Mn8@3247_g N_VSS_Mn8@3247_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3246 N_OUT8_Mn8@3246_d N_OUT7_Mn8@3246_g N_VSS_Mn8@3246_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3247 N_OUT8_Mp8@3247_d N_OUT7_Mp8@3247_g N_VDD_Mp8@3247_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3246 N_OUT8_Mp8@3246_d N_OUT7_Mp8@3246_g N_VDD_Mp8@3246_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3245 N_OUT8_Mn8@3245_d N_OUT7_Mn8@3245_g N_VSS_Mn8@3245_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3244 N_OUT8_Mn8@3244_d N_OUT7_Mn8@3244_g N_VSS_Mn8@3244_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3245 N_OUT8_Mp8@3245_d N_OUT7_Mp8@3245_g N_VDD_Mp8@3245_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3244 N_OUT8_Mp8@3244_d N_OUT7_Mp8@3244_g N_VDD_Mp8@3244_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3243 N_OUT8_Mn8@3243_d N_OUT7_Mn8@3243_g N_VSS_Mn8@3243_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3242 N_OUT8_Mn8@3242_d N_OUT7_Mn8@3242_g N_VSS_Mn8@3242_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3243 N_OUT8_Mp8@3243_d N_OUT7_Mp8@3243_g N_VDD_Mp8@3243_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3242 N_OUT8_Mp8@3242_d N_OUT7_Mp8@3242_g N_VDD_Mp8@3242_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3241 N_OUT8_Mn8@3241_d N_OUT7_Mn8@3241_g N_VSS_Mn8@3241_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3240 N_OUT8_Mn8@3240_d N_OUT7_Mn8@3240_g N_VSS_Mn8@3240_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3241 N_OUT8_Mp8@3241_d N_OUT7_Mp8@3241_g N_VDD_Mp8@3241_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3240 N_OUT8_Mp8@3240_d N_OUT7_Mp8@3240_g N_VDD_Mp8@3240_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3239 N_OUT8_Mn8@3239_d N_OUT7_Mn8@3239_g N_VSS_Mn8@3239_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3238 N_OUT8_Mn8@3238_d N_OUT7_Mn8@3238_g N_VSS_Mn8@3238_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3239 N_OUT8_Mp8@3239_d N_OUT7_Mp8@3239_g N_VDD_Mp8@3239_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3238 N_OUT8_Mp8@3238_d N_OUT7_Mp8@3238_g N_VDD_Mp8@3238_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3237 N_OUT8_Mn8@3237_d N_OUT7_Mn8@3237_g N_VSS_Mn8@3237_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3236 N_OUT8_Mn8@3236_d N_OUT7_Mn8@3236_g N_VSS_Mn8@3236_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3237 N_OUT8_Mp8@3237_d N_OUT7_Mp8@3237_g N_VDD_Mp8@3237_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3236 N_OUT8_Mp8@3236_d N_OUT7_Mp8@3236_g N_VDD_Mp8@3236_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3235 N_OUT8_Mn8@3235_d N_OUT7_Mn8@3235_g N_VSS_Mn8@3235_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3234 N_OUT8_Mn8@3234_d N_OUT7_Mn8@3234_g N_VSS_Mn8@3234_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3235 N_OUT8_Mp8@3235_d N_OUT7_Mp8@3235_g N_VDD_Mp8@3235_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3234 N_OUT8_Mp8@3234_d N_OUT7_Mp8@3234_g N_VDD_Mp8@3234_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3233 N_OUT8_Mn8@3233_d N_OUT7_Mn8@3233_g N_VSS_Mn8@3233_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3232 N_OUT8_Mn8@3232_d N_OUT7_Mn8@3232_g N_VSS_Mn8@3232_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3233 N_OUT8_Mp8@3233_d N_OUT7_Mp8@3233_g N_VDD_Mp8@3233_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3232 N_OUT8_Mp8@3232_d N_OUT7_Mp8@3232_g N_VDD_Mp8@3232_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3231 N_OUT8_Mn8@3231_d N_OUT7_Mn8@3231_g N_VSS_Mn8@3231_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3230 N_OUT8_Mn8@3230_d N_OUT7_Mn8@3230_g N_VSS_Mn8@3230_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3231 N_OUT8_Mp8@3231_d N_OUT7_Mp8@3231_g N_VDD_Mp8@3231_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3230 N_OUT8_Mp8@3230_d N_OUT7_Mp8@3230_g N_VDD_Mp8@3230_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3229 N_OUT8_Mn8@3229_d N_OUT7_Mn8@3229_g N_VSS_Mn8@3229_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3228 N_OUT8_Mn8@3228_d N_OUT7_Mn8@3228_g N_VSS_Mn8@3228_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3229 N_OUT8_Mp8@3229_d N_OUT7_Mp8@3229_g N_VDD_Mp8@3229_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3228 N_OUT8_Mp8@3228_d N_OUT7_Mp8@3228_g N_VDD_Mp8@3228_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3227 N_OUT8_Mn8@3227_d N_OUT7_Mn8@3227_g N_VSS_Mn8@3227_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3226 N_OUT8_Mn8@3226_d N_OUT7_Mn8@3226_g N_VSS_Mn8@3226_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3227 N_OUT8_Mp8@3227_d N_OUT7_Mp8@3227_g N_VDD_Mp8@3227_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3226 N_OUT8_Mp8@3226_d N_OUT7_Mp8@3226_g N_VDD_Mp8@3226_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3225 N_OUT8_Mn8@3225_d N_OUT7_Mn8@3225_g N_VSS_Mn8@3225_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3224 N_OUT8_Mn8@3224_d N_OUT7_Mn8@3224_g N_VSS_Mn8@3224_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3225 N_OUT8_Mp8@3225_d N_OUT7_Mp8@3225_g N_VDD_Mp8@3225_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3224 N_OUT8_Mp8@3224_d N_OUT7_Mp8@3224_g N_VDD_Mp8@3224_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3223 N_OUT8_Mn8@3223_d N_OUT7_Mn8@3223_g N_VSS_Mn8@3223_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3222 N_OUT8_Mn8@3222_d N_OUT7_Mn8@3222_g N_VSS_Mn8@3222_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3223 N_OUT8_Mp8@3223_d N_OUT7_Mp8@3223_g N_VDD_Mp8@3223_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3222 N_OUT8_Mp8@3222_d N_OUT7_Mp8@3222_g N_VDD_Mp8@3222_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3221 N_OUT8_Mn8@3221_d N_OUT7_Mn8@3221_g N_VSS_Mn8@3221_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3220 N_OUT8_Mn8@3220_d N_OUT7_Mn8@3220_g N_VSS_Mn8@3220_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3221 N_OUT8_Mp8@3221_d N_OUT7_Mp8@3221_g N_VDD_Mp8@3221_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3220 N_OUT8_Mp8@3220_d N_OUT7_Mp8@3220_g N_VDD_Mp8@3220_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3219 N_OUT8_Mn8@3219_d N_OUT7_Mn8@3219_g N_VSS_Mn8@3219_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3218 N_OUT8_Mn8@3218_d N_OUT7_Mn8@3218_g N_VSS_Mn8@3218_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3219 N_OUT8_Mp8@3219_d N_OUT7_Mp8@3219_g N_VDD_Mp8@3219_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3218 N_OUT8_Mp8@3218_d N_OUT7_Mp8@3218_g N_VDD_Mp8@3218_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3217 N_OUT8_Mn8@3217_d N_OUT7_Mn8@3217_g N_VSS_Mn8@3217_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3216 N_OUT8_Mn8@3216_d N_OUT7_Mn8@3216_g N_VSS_Mn8@3216_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3217 N_OUT8_Mp8@3217_d N_OUT7_Mp8@3217_g N_VDD_Mp8@3217_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3216 N_OUT8_Mp8@3216_d N_OUT7_Mp8@3216_g N_VDD_Mp8@3216_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3215 N_OUT8_Mn8@3215_d N_OUT7_Mn8@3215_g N_VSS_Mn8@3215_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3214 N_OUT8_Mn8@3214_d N_OUT7_Mn8@3214_g N_VSS_Mn8@3214_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3215 N_OUT8_Mp8@3215_d N_OUT7_Mp8@3215_g N_VDD_Mp8@3215_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3214 N_OUT8_Mp8@3214_d N_OUT7_Mp8@3214_g N_VDD_Mp8@3214_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3213 N_OUT8_Mn8@3213_d N_OUT7_Mn8@3213_g N_VSS_Mn8@3213_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3212 N_OUT8_Mn8@3212_d N_OUT7_Mn8@3212_g N_VSS_Mn8@3212_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3213 N_OUT8_Mp8@3213_d N_OUT7_Mp8@3213_g N_VDD_Mp8@3213_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3212 N_OUT8_Mp8@3212_d N_OUT7_Mp8@3212_g N_VDD_Mp8@3212_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3211 N_OUT8_Mn8@3211_d N_OUT7_Mn8@3211_g N_VSS_Mn8@3211_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3210 N_OUT8_Mn8@3210_d N_OUT7_Mn8@3210_g N_VSS_Mn8@3210_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3211 N_OUT8_Mp8@3211_d N_OUT7_Mp8@3211_g N_VDD_Mp8@3211_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3210 N_OUT8_Mp8@3210_d N_OUT7_Mp8@3210_g N_VDD_Mp8@3210_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3209 N_OUT8_Mn8@3209_d N_OUT7_Mn8@3209_g N_VSS_Mn8@3209_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3208 N_OUT8_Mn8@3208_d N_OUT7_Mn8@3208_g N_VSS_Mn8@3208_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3209 N_OUT8_Mp8@3209_d N_OUT7_Mp8@3209_g N_VDD_Mp8@3209_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3208 N_OUT8_Mp8@3208_d N_OUT7_Mp8@3208_g N_VDD_Mp8@3208_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3207 N_OUT8_Mn8@3207_d N_OUT7_Mn8@3207_g N_VSS_Mn8@3207_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3206 N_OUT8_Mn8@3206_d N_OUT7_Mn8@3206_g N_VSS_Mn8@3206_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3207 N_OUT8_Mp8@3207_d N_OUT7_Mp8@3207_g N_VDD_Mp8@3207_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3206 N_OUT8_Mp8@3206_d N_OUT7_Mp8@3206_g N_VDD_Mp8@3206_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3205 N_OUT8_Mn8@3205_d N_OUT7_Mn8@3205_g N_VSS_Mn8@3205_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3204 N_OUT8_Mn8@3204_d N_OUT7_Mn8@3204_g N_VSS_Mn8@3204_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3205 N_OUT8_Mp8@3205_d N_OUT7_Mp8@3205_g N_VDD_Mp8@3205_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3204 N_OUT8_Mp8@3204_d N_OUT7_Mp8@3204_g N_VDD_Mp8@3204_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3203 N_OUT8_Mn8@3203_d N_OUT7_Mn8@3203_g N_VSS_Mn8@3203_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3202 N_OUT8_Mn8@3202_d N_OUT7_Mn8@3202_g N_VSS_Mn8@3202_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3203 N_OUT8_Mp8@3203_d N_OUT7_Mp8@3203_g N_VDD_Mp8@3203_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3202 N_OUT8_Mp8@3202_d N_OUT7_Mp8@3202_g N_VDD_Mp8@3202_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3201 N_OUT8_Mn8@3201_d N_OUT7_Mn8@3201_g N_VSS_Mn8@3201_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3200 N_OUT8_Mn8@3200_d N_OUT7_Mn8@3200_g N_VSS_Mn8@3200_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3201 N_OUT8_Mp8@3201_d N_OUT7_Mp8@3201_g N_VDD_Mp8@3201_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3200 N_OUT8_Mp8@3200_d N_OUT7_Mp8@3200_g N_VDD_Mp8@3200_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3199 N_OUT8_Mn8@3199_d N_OUT7_Mn8@3199_g N_VSS_Mn8@3199_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3198 N_OUT8_Mn8@3198_d N_OUT7_Mn8@3198_g N_VSS_Mn8@3198_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3199 N_OUT8_Mp8@3199_d N_OUT7_Mp8@3199_g N_VDD_Mp8@3199_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3198 N_OUT8_Mp8@3198_d N_OUT7_Mp8@3198_g N_VDD_Mp8@3198_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3197 N_OUT8_Mn8@3197_d N_OUT7_Mn8@3197_g N_VSS_Mn8@3197_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3196 N_OUT8_Mn8@3196_d N_OUT7_Mn8@3196_g N_VSS_Mn8@3196_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3197 N_OUT8_Mp8@3197_d N_OUT7_Mp8@3197_g N_VDD_Mp8@3197_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3196 N_OUT8_Mp8@3196_d N_OUT7_Mp8@3196_g N_VDD_Mp8@3196_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3195 N_OUT8_Mn8@3195_d N_OUT7_Mn8@3195_g N_VSS_Mn8@3195_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3194 N_OUT8_Mn8@3194_d N_OUT7_Mn8@3194_g N_VSS_Mn8@3194_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3195 N_OUT8_Mp8@3195_d N_OUT7_Mp8@3195_g N_VDD_Mp8@3195_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3194 N_OUT8_Mp8@3194_d N_OUT7_Mp8@3194_g N_VDD_Mp8@3194_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3193 N_OUT8_Mn8@3193_d N_OUT7_Mn8@3193_g N_VSS_Mn8@3193_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3192 N_OUT8_Mn8@3192_d N_OUT7_Mn8@3192_g N_VSS_Mn8@3192_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3193 N_OUT8_Mp8@3193_d N_OUT7_Mp8@3193_g N_VDD_Mp8@3193_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3192 N_OUT8_Mp8@3192_d N_OUT7_Mp8@3192_g N_VDD_Mp8@3192_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3191 N_OUT8_Mn8@3191_d N_OUT7_Mn8@3191_g N_VSS_Mn8@3191_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3190 N_OUT8_Mn8@3190_d N_OUT7_Mn8@3190_g N_VSS_Mn8@3190_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3191 N_OUT8_Mp8@3191_d N_OUT7_Mp8@3191_g N_VDD_Mp8@3191_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3190 N_OUT8_Mp8@3190_d N_OUT7_Mp8@3190_g N_VDD_Mp8@3190_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3189 N_OUT8_Mn8@3189_d N_OUT7_Mn8@3189_g N_VSS_Mn8@3189_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3188 N_OUT8_Mn8@3188_d N_OUT7_Mn8@3188_g N_VSS_Mn8@3188_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3189 N_OUT8_Mp8@3189_d N_OUT7_Mp8@3189_g N_VDD_Mp8@3189_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3188 N_OUT8_Mp8@3188_d N_OUT7_Mp8@3188_g N_VDD_Mp8@3188_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3187 N_OUT8_Mn8@3187_d N_OUT7_Mn8@3187_g N_VSS_Mn8@3187_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3186 N_OUT8_Mn8@3186_d N_OUT7_Mn8@3186_g N_VSS_Mn8@3186_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3187 N_OUT8_Mp8@3187_d N_OUT7_Mp8@3187_g N_VDD_Mp8@3187_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3186 N_OUT8_Mp8@3186_d N_OUT7_Mp8@3186_g N_VDD_Mp8@3186_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3185 N_OUT8_Mn8@3185_d N_OUT7_Mn8@3185_g N_VSS_Mn8@3185_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3184 N_OUT8_Mn8@3184_d N_OUT7_Mn8@3184_g N_VSS_Mn8@3184_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3185 N_OUT8_Mp8@3185_d N_OUT7_Mp8@3185_g N_VDD_Mp8@3185_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3184 N_OUT8_Mp8@3184_d N_OUT7_Mp8@3184_g N_VDD_Mp8@3184_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3183 N_OUT8_Mn8@3183_d N_OUT7_Mn8@3183_g N_VSS_Mn8@3183_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3182 N_OUT8_Mn8@3182_d N_OUT7_Mn8@3182_g N_VSS_Mn8@3182_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3183 N_OUT8_Mp8@3183_d N_OUT7_Mp8@3183_g N_VDD_Mp8@3183_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3182 N_OUT8_Mp8@3182_d N_OUT7_Mp8@3182_g N_VDD_Mp8@3182_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3181 N_OUT8_Mn8@3181_d N_OUT7_Mn8@3181_g N_VSS_Mn8@3181_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3180 N_OUT8_Mn8@3180_d N_OUT7_Mn8@3180_g N_VSS_Mn8@3180_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3181 N_OUT8_Mp8@3181_d N_OUT7_Mp8@3181_g N_VDD_Mp8@3181_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3180 N_OUT8_Mp8@3180_d N_OUT7_Mp8@3180_g N_VDD_Mp8@3180_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3179 N_OUT8_Mn8@3179_d N_OUT7_Mn8@3179_g N_VSS_Mn8@3179_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3178 N_OUT8_Mn8@3178_d N_OUT7_Mn8@3178_g N_VSS_Mn8@3178_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3179 N_OUT8_Mp8@3179_d N_OUT7_Mp8@3179_g N_VDD_Mp8@3179_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3178 N_OUT8_Mp8@3178_d N_OUT7_Mp8@3178_g N_VDD_Mp8@3178_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3177 N_OUT8_Mn8@3177_d N_OUT7_Mn8@3177_g N_VSS_Mn8@3177_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3176 N_OUT8_Mn8@3176_d N_OUT7_Mn8@3176_g N_VSS_Mn8@3176_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3177 N_OUT8_Mp8@3177_d N_OUT7_Mp8@3177_g N_VDD_Mp8@3177_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3176 N_OUT8_Mp8@3176_d N_OUT7_Mp8@3176_g N_VDD_Mp8@3176_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3175 N_OUT8_Mn8@3175_d N_OUT7_Mn8@3175_g N_VSS_Mn8@3175_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3174 N_OUT8_Mn8@3174_d N_OUT7_Mn8@3174_g N_VSS_Mn8@3174_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3175 N_OUT8_Mp8@3175_d N_OUT7_Mp8@3175_g N_VDD_Mp8@3175_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3174 N_OUT8_Mp8@3174_d N_OUT7_Mp8@3174_g N_VDD_Mp8@3174_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3173 N_OUT8_Mn8@3173_d N_OUT7_Mn8@3173_g N_VSS_Mn8@3173_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3172 N_OUT8_Mn8@3172_d N_OUT7_Mn8@3172_g N_VSS_Mn8@3172_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3173 N_OUT8_Mp8@3173_d N_OUT7_Mp8@3173_g N_VDD_Mp8@3173_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3172 N_OUT8_Mp8@3172_d N_OUT7_Mp8@3172_g N_VDD_Mp8@3172_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3171 N_OUT8_Mn8@3171_d N_OUT7_Mn8@3171_g N_VSS_Mn8@3171_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3170 N_OUT8_Mn8@3170_d N_OUT7_Mn8@3170_g N_VSS_Mn8@3170_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3171 N_OUT8_Mp8@3171_d N_OUT7_Mp8@3171_g N_VDD_Mp8@3171_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3170 N_OUT8_Mp8@3170_d N_OUT7_Mp8@3170_g N_VDD_Mp8@3170_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3169 N_OUT8_Mn8@3169_d N_OUT7_Mn8@3169_g N_VSS_Mn8@3169_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3168 N_OUT8_Mn8@3168_d N_OUT7_Mn8@3168_g N_VSS_Mn8@3168_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3169 N_OUT8_Mp8@3169_d N_OUT7_Mp8@3169_g N_VDD_Mp8@3169_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3168 N_OUT8_Mp8@3168_d N_OUT7_Mp8@3168_g N_VDD_Mp8@3168_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3167 N_OUT8_Mn8@3167_d N_OUT7_Mn8@3167_g N_VSS_Mn8@3167_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3166 N_OUT8_Mn8@3166_d N_OUT7_Mn8@3166_g N_VSS_Mn8@3166_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3167 N_OUT8_Mp8@3167_d N_OUT7_Mp8@3167_g N_VDD_Mp8@3167_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3166 N_OUT8_Mp8@3166_d N_OUT7_Mp8@3166_g N_VDD_Mp8@3166_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3165 N_OUT8_Mn8@3165_d N_OUT7_Mn8@3165_g N_VSS_Mn8@3165_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3164 N_OUT8_Mn8@3164_d N_OUT7_Mn8@3164_g N_VSS_Mn8@3164_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3165 N_OUT8_Mp8@3165_d N_OUT7_Mp8@3165_g N_VDD_Mp8@3165_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3164 N_OUT8_Mp8@3164_d N_OUT7_Mp8@3164_g N_VDD_Mp8@3164_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3163 N_OUT8_Mn8@3163_d N_OUT7_Mn8@3163_g N_VSS_Mn8@3163_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3162 N_OUT8_Mn8@3162_d N_OUT7_Mn8@3162_g N_VSS_Mn8@3162_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3163 N_OUT8_Mp8@3163_d N_OUT7_Mp8@3163_g N_VDD_Mp8@3163_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3162 N_OUT8_Mp8@3162_d N_OUT7_Mp8@3162_g N_VDD_Mp8@3162_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3161 N_OUT8_Mn8@3161_d N_OUT7_Mn8@3161_g N_VSS_Mn8@3161_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3160 N_OUT8_Mn8@3160_d N_OUT7_Mn8@3160_g N_VSS_Mn8@3160_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3161 N_OUT8_Mp8@3161_d N_OUT7_Mp8@3161_g N_VDD_Mp8@3161_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3160 N_OUT8_Mp8@3160_d N_OUT7_Mp8@3160_g N_VDD_Mp8@3160_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3159 N_OUT8_Mn8@3159_d N_OUT7_Mn8@3159_g N_VSS_Mn8@3159_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3158 N_OUT8_Mn8@3158_d N_OUT7_Mn8@3158_g N_VSS_Mn8@3158_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3159 N_OUT8_Mp8@3159_d N_OUT7_Mp8@3159_g N_VDD_Mp8@3159_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3158 N_OUT8_Mp8@3158_d N_OUT7_Mp8@3158_g N_VDD_Mp8@3158_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3157 N_OUT8_Mn8@3157_d N_OUT7_Mn8@3157_g N_VSS_Mn8@3157_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3156 N_OUT8_Mn8@3156_d N_OUT7_Mn8@3156_g N_VSS_Mn8@3156_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3157 N_OUT8_Mp8@3157_d N_OUT7_Mp8@3157_g N_VDD_Mp8@3157_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3156 N_OUT8_Mp8@3156_d N_OUT7_Mp8@3156_g N_VDD_Mp8@3156_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3155 N_OUT8_Mn8@3155_d N_OUT7_Mn8@3155_g N_VSS_Mn8@3155_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3154 N_OUT8_Mn8@3154_d N_OUT7_Mn8@3154_g N_VSS_Mn8@3154_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3155 N_OUT8_Mp8@3155_d N_OUT7_Mp8@3155_g N_VDD_Mp8@3155_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3154 N_OUT8_Mp8@3154_d N_OUT7_Mp8@3154_g N_VDD_Mp8@3154_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3153 N_OUT8_Mn8@3153_d N_OUT7_Mn8@3153_g N_VSS_Mn8@3153_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3152 N_OUT8_Mn8@3152_d N_OUT7_Mn8@3152_g N_VSS_Mn8@3152_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3153 N_OUT8_Mp8@3153_d N_OUT7_Mp8@3153_g N_VDD_Mp8@3153_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3152 N_OUT8_Mp8@3152_d N_OUT7_Mp8@3152_g N_VDD_Mp8@3152_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3151 N_OUT8_Mn8@3151_d N_OUT7_Mn8@3151_g N_VSS_Mn8@3151_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3150 N_OUT8_Mn8@3150_d N_OUT7_Mn8@3150_g N_VSS_Mn8@3150_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3151 N_OUT8_Mp8@3151_d N_OUT7_Mp8@3151_g N_VDD_Mp8@3151_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3150 N_OUT8_Mp8@3150_d N_OUT7_Mp8@3150_g N_VDD_Mp8@3150_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3149 N_OUT8_Mn8@3149_d N_OUT7_Mn8@3149_g N_VSS_Mn8@3149_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3148 N_OUT8_Mn8@3148_d N_OUT7_Mn8@3148_g N_VSS_Mn8@3148_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3149 N_OUT8_Mp8@3149_d N_OUT7_Mp8@3149_g N_VDD_Mp8@3149_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3148 N_OUT8_Mp8@3148_d N_OUT7_Mp8@3148_g N_VDD_Mp8@3148_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3147 N_OUT8_Mn8@3147_d N_OUT7_Mn8@3147_g N_VSS_Mn8@3147_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3146 N_OUT8_Mn8@3146_d N_OUT7_Mn8@3146_g N_VSS_Mn8@3146_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3147 N_OUT8_Mp8@3147_d N_OUT7_Mp8@3147_g N_VDD_Mp8@3147_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3146 N_OUT8_Mp8@3146_d N_OUT7_Mp8@3146_g N_VDD_Mp8@3146_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3145 N_OUT8_Mn8@3145_d N_OUT7_Mn8@3145_g N_VSS_Mn8@3145_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3144 N_OUT8_Mn8@3144_d N_OUT7_Mn8@3144_g N_VSS_Mn8@3144_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3145 N_OUT8_Mp8@3145_d N_OUT7_Mp8@3145_g N_VDD_Mp8@3145_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3144 N_OUT8_Mp8@3144_d N_OUT7_Mp8@3144_g N_VDD_Mp8@3144_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3143 N_OUT8_Mn8@3143_d N_OUT7_Mn8@3143_g N_VSS_Mn8@3143_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3142 N_OUT8_Mn8@3142_d N_OUT7_Mn8@3142_g N_VSS_Mn8@3142_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3143 N_OUT8_Mp8@3143_d N_OUT7_Mp8@3143_g N_VDD_Mp8@3143_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3142 N_OUT8_Mp8@3142_d N_OUT7_Mp8@3142_g N_VDD_Mp8@3142_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3141 N_OUT8_Mn8@3141_d N_OUT7_Mn8@3141_g N_VSS_Mn8@3141_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3140 N_OUT8_Mn8@3140_d N_OUT7_Mn8@3140_g N_VSS_Mn8@3140_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3141 N_OUT8_Mp8@3141_d N_OUT7_Mp8@3141_g N_VDD_Mp8@3141_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3140 N_OUT8_Mp8@3140_d N_OUT7_Mp8@3140_g N_VDD_Mp8@3140_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3139 N_OUT8_Mn8@3139_d N_OUT7_Mn8@3139_g N_VSS_Mn8@3139_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3138 N_OUT8_Mn8@3138_d N_OUT7_Mn8@3138_g N_VSS_Mn8@3138_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3139 N_OUT8_Mp8@3139_d N_OUT7_Mp8@3139_g N_VDD_Mp8@3139_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3138 N_OUT8_Mp8@3138_d N_OUT7_Mp8@3138_g N_VDD_Mp8@3138_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3137 N_OUT8_Mn8@3137_d N_OUT7_Mn8@3137_g N_VSS_Mn8@3137_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3136 N_OUT8_Mn8@3136_d N_OUT7_Mn8@3136_g N_VSS_Mn8@3136_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3137 N_OUT8_Mp8@3137_d N_OUT7_Mp8@3137_g N_VDD_Mp8@3137_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3136 N_OUT8_Mp8@3136_d N_OUT7_Mp8@3136_g N_VDD_Mp8@3136_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3135 N_OUT8_Mn8@3135_d N_OUT7_Mn8@3135_g N_VSS_Mn8@3135_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3134 N_OUT8_Mn8@3134_d N_OUT7_Mn8@3134_g N_VSS_Mn8@3134_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3135 N_OUT8_Mp8@3135_d N_OUT7_Mp8@3135_g N_VDD_Mp8@3135_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3134 N_OUT8_Mp8@3134_d N_OUT7_Mp8@3134_g N_VDD_Mp8@3134_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3133 N_OUT8_Mn8@3133_d N_OUT7_Mn8@3133_g N_VSS_Mn8@3133_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3132 N_OUT8_Mn8@3132_d N_OUT7_Mn8@3132_g N_VSS_Mn8@3132_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3133 N_OUT8_Mp8@3133_d N_OUT7_Mp8@3133_g N_VDD_Mp8@3133_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3132 N_OUT8_Mp8@3132_d N_OUT7_Mp8@3132_g N_VDD_Mp8@3132_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3131 N_OUT8_Mn8@3131_d N_OUT7_Mn8@3131_g N_VSS_Mn8@3131_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3130 N_OUT8_Mn8@3130_d N_OUT7_Mn8@3130_g N_VSS_Mn8@3130_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3131 N_OUT8_Mp8@3131_d N_OUT7_Mp8@3131_g N_VDD_Mp8@3131_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3130 N_OUT8_Mp8@3130_d N_OUT7_Mp8@3130_g N_VDD_Mp8@3130_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3129 N_OUT8_Mn8@3129_d N_OUT7_Mn8@3129_g N_VSS_Mn8@3129_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3128 N_OUT8_Mn8@3128_d N_OUT7_Mn8@3128_g N_VSS_Mn8@3128_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3129 N_OUT8_Mp8@3129_d N_OUT7_Mp8@3129_g N_VDD_Mp8@3129_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3128 N_OUT8_Mp8@3128_d N_OUT7_Mp8@3128_g N_VDD_Mp8@3128_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3127 N_OUT8_Mn8@3127_d N_OUT7_Mn8@3127_g N_VSS_Mn8@3127_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3126 N_OUT8_Mn8@3126_d N_OUT7_Mn8@3126_g N_VSS_Mn8@3126_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3127 N_OUT8_Mp8@3127_d N_OUT7_Mp8@3127_g N_VDD_Mp8@3127_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3126 N_OUT8_Mp8@3126_d N_OUT7_Mp8@3126_g N_VDD_Mp8@3126_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3125 N_OUT8_Mn8@3125_d N_OUT7_Mn8@3125_g N_VSS_Mn8@3125_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3124 N_OUT8_Mn8@3124_d N_OUT7_Mn8@3124_g N_VSS_Mn8@3124_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3125 N_OUT8_Mp8@3125_d N_OUT7_Mp8@3125_g N_VDD_Mp8@3125_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3124 N_OUT8_Mp8@3124_d N_OUT7_Mp8@3124_g N_VDD_Mp8@3124_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3123 N_OUT8_Mn8@3123_d N_OUT7_Mn8@3123_g N_VSS_Mn8@3123_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3122 N_OUT8_Mn8@3122_d N_OUT7_Mn8@3122_g N_VSS_Mn8@3122_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3123 N_OUT8_Mp8@3123_d N_OUT7_Mp8@3123_g N_VDD_Mp8@3123_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3122 N_OUT8_Mp8@3122_d N_OUT7_Mp8@3122_g N_VDD_Mp8@3122_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3121 N_OUT8_Mn8@3121_d N_OUT7_Mn8@3121_g N_VSS_Mn8@3121_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3120 N_OUT8_Mn8@3120_d N_OUT7_Mn8@3120_g N_VSS_Mn8@3120_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3121 N_OUT8_Mp8@3121_d N_OUT7_Mp8@3121_g N_VDD_Mp8@3121_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3120 N_OUT8_Mp8@3120_d N_OUT7_Mp8@3120_g N_VDD_Mp8@3120_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3119 N_OUT8_Mn8@3119_d N_OUT7_Mn8@3119_g N_VSS_Mn8@3119_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3118 N_OUT8_Mn8@3118_d N_OUT7_Mn8@3118_g N_VSS_Mn8@3118_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3119 N_OUT8_Mp8@3119_d N_OUT7_Mp8@3119_g N_VDD_Mp8@3119_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3118 N_OUT8_Mp8@3118_d N_OUT7_Mp8@3118_g N_VDD_Mp8@3118_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3117 N_OUT8_Mn8@3117_d N_OUT7_Mn8@3117_g N_VSS_Mn8@3117_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3116 N_OUT8_Mn8@3116_d N_OUT7_Mn8@3116_g N_VSS_Mn8@3116_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3117 N_OUT8_Mp8@3117_d N_OUT7_Mp8@3117_g N_VDD_Mp8@3117_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3116 N_OUT8_Mp8@3116_d N_OUT7_Mp8@3116_g N_VDD_Mp8@3116_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3115 N_OUT8_Mn8@3115_d N_OUT7_Mn8@3115_g N_VSS_Mn8@3115_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3114 N_OUT8_Mn8@3114_d N_OUT7_Mn8@3114_g N_VSS_Mn8@3114_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3115 N_OUT8_Mp8@3115_d N_OUT7_Mp8@3115_g N_VDD_Mp8@3115_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3114 N_OUT8_Mp8@3114_d N_OUT7_Mp8@3114_g N_VDD_Mp8@3114_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3113 N_OUT8_Mn8@3113_d N_OUT7_Mn8@3113_g N_VSS_Mn8@3113_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3112 N_OUT8_Mn8@3112_d N_OUT7_Mn8@3112_g N_VSS_Mn8@3112_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3113 N_OUT8_Mp8@3113_d N_OUT7_Mp8@3113_g N_VDD_Mp8@3113_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3112 N_OUT8_Mp8@3112_d N_OUT7_Mp8@3112_g N_VDD_Mp8@3112_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3111 N_OUT8_Mn8@3111_d N_OUT7_Mn8@3111_g N_VSS_Mn8@3111_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3110 N_OUT8_Mn8@3110_d N_OUT7_Mn8@3110_g N_VSS_Mn8@3110_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3111 N_OUT8_Mp8@3111_d N_OUT7_Mp8@3111_g N_VDD_Mp8@3111_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3110 N_OUT8_Mp8@3110_d N_OUT7_Mp8@3110_g N_VDD_Mp8@3110_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3109 N_OUT8_Mn8@3109_d N_OUT7_Mn8@3109_g N_VSS_Mn8@3109_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3108 N_OUT8_Mn8@3108_d N_OUT7_Mn8@3108_g N_VSS_Mn8@3108_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3109 N_OUT8_Mp8@3109_d N_OUT7_Mp8@3109_g N_VDD_Mp8@3109_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3108 N_OUT8_Mp8@3108_d N_OUT7_Mp8@3108_g N_VDD_Mp8@3108_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3107 N_OUT8_Mn8@3107_d N_OUT7_Mn8@3107_g N_VSS_Mn8@3107_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3106 N_OUT8_Mn8@3106_d N_OUT7_Mn8@3106_g N_VSS_Mn8@3106_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3107 N_OUT8_Mp8@3107_d N_OUT7_Mp8@3107_g N_VDD_Mp8@3107_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3106 N_OUT8_Mp8@3106_d N_OUT7_Mp8@3106_g N_VDD_Mp8@3106_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3105 N_OUT8_Mn8@3105_d N_OUT7_Mn8@3105_g N_VSS_Mn8@3105_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3104 N_OUT8_Mn8@3104_d N_OUT7_Mn8@3104_g N_VSS_Mn8@3104_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3105 N_OUT8_Mp8@3105_d N_OUT7_Mp8@3105_g N_VDD_Mp8@3105_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3104 N_OUT8_Mp8@3104_d N_OUT7_Mp8@3104_g N_VDD_Mp8@3104_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3103 N_OUT8_Mn8@3103_d N_OUT7_Mn8@3103_g N_VSS_Mn8@3103_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3102 N_OUT8_Mn8@3102_d N_OUT7_Mn8@3102_g N_VSS_Mn8@3102_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3103 N_OUT8_Mp8@3103_d N_OUT7_Mp8@3103_g N_VDD_Mp8@3103_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3102 N_OUT8_Mp8@3102_d N_OUT7_Mp8@3102_g N_VDD_Mp8@3102_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3101 N_OUT8_Mn8@3101_d N_OUT7_Mn8@3101_g N_VSS_Mn8@3101_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3100 N_OUT8_Mn8@3100_d N_OUT7_Mn8@3100_g N_VSS_Mn8@3100_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3101 N_OUT8_Mp8@3101_d N_OUT7_Mp8@3101_g N_VDD_Mp8@3101_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3100 N_OUT8_Mp8@3100_d N_OUT7_Mp8@3100_g N_VDD_Mp8@3100_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3099 N_OUT8_Mn8@3099_d N_OUT7_Mn8@3099_g N_VSS_Mn8@3099_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3098 N_OUT8_Mn8@3098_d N_OUT7_Mn8@3098_g N_VSS_Mn8@3098_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3099 N_OUT8_Mp8@3099_d N_OUT7_Mp8@3099_g N_VDD_Mp8@3099_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3098 N_OUT8_Mp8@3098_d N_OUT7_Mp8@3098_g N_VDD_Mp8@3098_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3097 N_OUT8_Mn8@3097_d N_OUT7_Mn8@3097_g N_VSS_Mn8@3097_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3096 N_OUT8_Mn8@3096_d N_OUT7_Mn8@3096_g N_VSS_Mn8@3096_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3097 N_OUT8_Mp8@3097_d N_OUT7_Mp8@3097_g N_VDD_Mp8@3097_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3096 N_OUT8_Mp8@3096_d N_OUT7_Mp8@3096_g N_VDD_Mp8@3096_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3095 N_OUT8_Mn8@3095_d N_OUT7_Mn8@3095_g N_VSS_Mn8@3095_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3094 N_OUT8_Mn8@3094_d N_OUT7_Mn8@3094_g N_VSS_Mn8@3094_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3095 N_OUT8_Mp8@3095_d N_OUT7_Mp8@3095_g N_VDD_Mp8@3095_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3094 N_OUT8_Mp8@3094_d N_OUT7_Mp8@3094_g N_VDD_Mp8@3094_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3093 N_OUT8_Mn8@3093_d N_OUT7_Mn8@3093_g N_VSS_Mn8@3093_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3092 N_OUT8_Mn8@3092_d N_OUT7_Mn8@3092_g N_VSS_Mn8@3092_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3093 N_OUT8_Mp8@3093_d N_OUT7_Mp8@3093_g N_VDD_Mp8@3093_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3092 N_OUT8_Mp8@3092_d N_OUT7_Mp8@3092_g N_VDD_Mp8@3092_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3091 N_OUT8_Mn8@3091_d N_OUT7_Mn8@3091_g N_VSS_Mn8@3091_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3090 N_OUT8_Mn8@3090_d N_OUT7_Mn8@3090_g N_VSS_Mn8@3090_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3091 N_OUT8_Mp8@3091_d N_OUT7_Mp8@3091_g N_VDD_Mp8@3091_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3090 N_OUT8_Mp8@3090_d N_OUT7_Mp8@3090_g N_VDD_Mp8@3090_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3089 N_OUT8_Mn8@3089_d N_OUT7_Mn8@3089_g N_VSS_Mn8@3089_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3088 N_OUT8_Mn8@3088_d N_OUT7_Mn8@3088_g N_VSS_Mn8@3088_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3089 N_OUT8_Mp8@3089_d N_OUT7_Mp8@3089_g N_VDD_Mp8@3089_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3088 N_OUT8_Mp8@3088_d N_OUT7_Mp8@3088_g N_VDD_Mp8@3088_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3087 N_OUT8_Mn8@3087_d N_OUT7_Mn8@3087_g N_VSS_Mn8@3087_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3086 N_OUT8_Mn8@3086_d N_OUT7_Mn8@3086_g N_VSS_Mn8@3086_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3087 N_OUT8_Mp8@3087_d N_OUT7_Mp8@3087_g N_VDD_Mp8@3087_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3086 N_OUT8_Mp8@3086_d N_OUT7_Mp8@3086_g N_VDD_Mp8@3086_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3085 N_OUT8_Mn8@3085_d N_OUT7_Mn8@3085_g N_VSS_Mn8@3085_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3084 N_OUT8_Mn8@3084_d N_OUT7_Mn8@3084_g N_VSS_Mn8@3084_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3085 N_OUT8_Mp8@3085_d N_OUT7_Mp8@3085_g N_VDD_Mp8@3085_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3084 N_OUT8_Mp8@3084_d N_OUT7_Mp8@3084_g N_VDD_Mp8@3084_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3083 N_OUT8_Mn8@3083_d N_OUT7_Mn8@3083_g N_VSS_Mn8@3083_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3082 N_OUT8_Mn8@3082_d N_OUT7_Mn8@3082_g N_VSS_Mn8@3082_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3083 N_OUT8_Mp8@3083_d N_OUT7_Mp8@3083_g N_VDD_Mp8@3083_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3082 N_OUT8_Mp8@3082_d N_OUT7_Mp8@3082_g N_VDD_Mp8@3082_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3081 N_OUT8_Mn8@3081_d N_OUT7_Mn8@3081_g N_VSS_Mn8@3081_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3080 N_OUT8_Mn8@3080_d N_OUT7_Mn8@3080_g N_VSS_Mn8@3080_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3081 N_OUT8_Mp8@3081_d N_OUT7_Mp8@3081_g N_VDD_Mp8@3081_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3080 N_OUT8_Mp8@3080_d N_OUT7_Mp8@3080_g N_VDD_Mp8@3080_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3079 N_OUT8_Mn8@3079_d N_OUT7_Mn8@3079_g N_VSS_Mn8@3079_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3078 N_OUT8_Mn8@3078_d N_OUT7_Mn8@3078_g N_VSS_Mn8@3078_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3079 N_OUT8_Mp8@3079_d N_OUT7_Mp8@3079_g N_VDD_Mp8@3079_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3078 N_OUT8_Mp8@3078_d N_OUT7_Mp8@3078_g N_VDD_Mp8@3078_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3077 N_OUT8_Mn8@3077_d N_OUT7_Mn8@3077_g N_VSS_Mn8@3077_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3076 N_OUT8_Mn8@3076_d N_OUT7_Mn8@3076_g N_VSS_Mn8@3076_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3077 N_OUT8_Mp8@3077_d N_OUT7_Mp8@3077_g N_VDD_Mp8@3077_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3076 N_OUT8_Mp8@3076_d N_OUT7_Mp8@3076_g N_VDD_Mp8@3076_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3075 N_OUT8_Mn8@3075_d N_OUT7_Mn8@3075_g N_VSS_Mn8@3075_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3074 N_OUT8_Mn8@3074_d N_OUT7_Mn8@3074_g N_VSS_Mn8@3074_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3075 N_OUT8_Mp8@3075_d N_OUT7_Mp8@3075_g N_VDD_Mp8@3075_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3074 N_OUT8_Mp8@3074_d N_OUT7_Mp8@3074_g N_VDD_Mp8@3074_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4609 N_OUT9_Mn9@4609_d N_OUT8_Mn9@4609_g N_VSS_Mn9@4609_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4608 N_OUT9_Mn9@4608_d N_OUT8_Mn9@4608_g N_VSS_Mn9@4608_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4609 N_OUT9_Mp9@4609_d N_OUT8_Mp9@4609_g N_VDD_Mp9@4609_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4608 N_OUT9_Mp9@4608_d N_OUT8_Mp9@4608_g N_VDD_Mp9@4608_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4607 N_OUT9_Mn9@4607_d N_OUT8_Mn9@4607_g N_VSS_Mn9@4607_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4606 N_OUT9_Mn9@4606_d N_OUT8_Mn9@4606_g N_VSS_Mn9@4606_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4607 N_OUT9_Mp9@4607_d N_OUT8_Mp9@4607_g N_VDD_Mp9@4607_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4606 N_OUT9_Mp9@4606_d N_OUT8_Mp9@4606_g N_VDD_Mp9@4606_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4605 N_OUT9_Mn9@4605_d N_OUT8_Mn9@4605_g N_VSS_Mn9@4605_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4604 N_OUT9_Mn9@4604_d N_OUT8_Mn9@4604_g N_VSS_Mn9@4604_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4605 N_OUT9_Mp9@4605_d N_OUT8_Mp9@4605_g N_VDD_Mp9@4605_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4604 N_OUT9_Mp9@4604_d N_OUT8_Mp9@4604_g N_VDD_Mp9@4604_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4603 N_OUT9_Mn9@4603_d N_OUT8_Mn9@4603_g N_VSS_Mn9@4603_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4602 N_OUT9_Mn9@4602_d N_OUT8_Mn9@4602_g N_VSS_Mn9@4602_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4603 N_OUT9_Mp9@4603_d N_OUT8_Mp9@4603_g N_VDD_Mp9@4603_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4602 N_OUT9_Mp9@4602_d N_OUT8_Mp9@4602_g N_VDD_Mp9@4602_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4601 N_OUT9_Mn9@4601_d N_OUT8_Mn9@4601_g N_VSS_Mn9@4601_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4600 N_OUT9_Mn9@4600_d N_OUT8_Mn9@4600_g N_VSS_Mn9@4600_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4601 N_OUT9_Mp9@4601_d N_OUT8_Mp9@4601_g N_VDD_Mp9@4601_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4600 N_OUT9_Mp9@4600_d N_OUT8_Mp9@4600_g N_VDD_Mp9@4600_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4599 N_OUT9_Mn9@4599_d N_OUT8_Mn9@4599_g N_VSS_Mn9@4599_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4598 N_OUT9_Mn9@4598_d N_OUT8_Mn9@4598_g N_VSS_Mn9@4598_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4599 N_OUT9_Mp9@4599_d N_OUT8_Mp9@4599_g N_VDD_Mp9@4599_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4598 N_OUT9_Mp9@4598_d N_OUT8_Mp9@4598_g N_VDD_Mp9@4598_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4597 N_OUT9_Mn9@4597_d N_OUT8_Mn9@4597_g N_VSS_Mn9@4597_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4596 N_OUT9_Mn9@4596_d N_OUT8_Mn9@4596_g N_VSS_Mn9@4596_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4597 N_OUT9_Mp9@4597_d N_OUT8_Mp9@4597_g N_VDD_Mp9@4597_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4596 N_OUT9_Mp9@4596_d N_OUT8_Mp9@4596_g N_VDD_Mp9@4596_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4595 N_OUT9_Mn9@4595_d N_OUT8_Mn9@4595_g N_VSS_Mn9@4595_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4594 N_OUT9_Mn9@4594_d N_OUT8_Mn9@4594_g N_VSS_Mn9@4594_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4595 N_OUT9_Mp9@4595_d N_OUT8_Mp9@4595_g N_VDD_Mp9@4595_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4594 N_OUT9_Mp9@4594_d N_OUT8_Mp9@4594_g N_VDD_Mp9@4594_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4593 N_OUT9_Mn9@4593_d N_OUT8_Mn9@4593_g N_VSS_Mn9@4593_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4592 N_OUT9_Mn9@4592_d N_OUT8_Mn9@4592_g N_VSS_Mn9@4592_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4593 N_OUT9_Mp9@4593_d N_OUT8_Mp9@4593_g N_VDD_Mp9@4593_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4592 N_OUT9_Mp9@4592_d N_OUT8_Mp9@4592_g N_VDD_Mp9@4592_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4591 N_OUT9_Mn9@4591_d N_OUT8_Mn9@4591_g N_VSS_Mn9@4591_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4590 N_OUT9_Mn9@4590_d N_OUT8_Mn9@4590_g N_VSS_Mn9@4590_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4591 N_OUT9_Mp9@4591_d N_OUT8_Mp9@4591_g N_VDD_Mp9@4591_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4590 N_OUT9_Mp9@4590_d N_OUT8_Mp9@4590_g N_VDD_Mp9@4590_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4589 N_OUT9_Mn9@4589_d N_OUT8_Mn9@4589_g N_VSS_Mn9@4589_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4588 N_OUT9_Mn9@4588_d N_OUT8_Mn9@4588_g N_VSS_Mn9@4588_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4589 N_OUT9_Mp9@4589_d N_OUT8_Mp9@4589_g N_VDD_Mp9@4589_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4588 N_OUT9_Mp9@4588_d N_OUT8_Mp9@4588_g N_VDD_Mp9@4588_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4587 N_OUT9_Mn9@4587_d N_OUT8_Mn9@4587_g N_VSS_Mn9@4587_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4586 N_OUT9_Mn9@4586_d N_OUT8_Mn9@4586_g N_VSS_Mn9@4586_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4587 N_OUT9_Mp9@4587_d N_OUT8_Mp9@4587_g N_VDD_Mp9@4587_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4586 N_OUT9_Mp9@4586_d N_OUT8_Mp9@4586_g N_VDD_Mp9@4586_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4585 N_OUT9_Mn9@4585_d N_OUT8_Mn9@4585_g N_VSS_Mn9@4585_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4584 N_OUT9_Mn9@4584_d N_OUT8_Mn9@4584_g N_VSS_Mn9@4584_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4585 N_OUT9_Mp9@4585_d N_OUT8_Mp9@4585_g N_VDD_Mp9@4585_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4584 N_OUT9_Mp9@4584_d N_OUT8_Mp9@4584_g N_VDD_Mp9@4584_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4583 N_OUT9_Mn9@4583_d N_OUT8_Mn9@4583_g N_VSS_Mn9@4583_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4582 N_OUT9_Mn9@4582_d N_OUT8_Mn9@4582_g N_VSS_Mn9@4582_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4583 N_OUT9_Mp9@4583_d N_OUT8_Mp9@4583_g N_VDD_Mp9@4583_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4582 N_OUT9_Mp9@4582_d N_OUT8_Mp9@4582_g N_VDD_Mp9@4582_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4581 N_OUT9_Mn9@4581_d N_OUT8_Mn9@4581_g N_VSS_Mn9@4581_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4580 N_OUT9_Mn9@4580_d N_OUT8_Mn9@4580_g N_VSS_Mn9@4580_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4581 N_OUT9_Mp9@4581_d N_OUT8_Mp9@4581_g N_VDD_Mp9@4581_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4580 N_OUT9_Mp9@4580_d N_OUT8_Mp9@4580_g N_VDD_Mp9@4580_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4579 N_OUT9_Mn9@4579_d N_OUT8_Mn9@4579_g N_VSS_Mn9@4579_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4578 N_OUT9_Mn9@4578_d N_OUT8_Mn9@4578_g N_VSS_Mn9@4578_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4579 N_OUT9_Mp9@4579_d N_OUT8_Mp9@4579_g N_VDD_Mp9@4579_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4578 N_OUT9_Mp9@4578_d N_OUT8_Mp9@4578_g N_VDD_Mp9@4578_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4577 N_OUT9_Mn9@4577_d N_OUT8_Mn9@4577_g N_VSS_Mn9@4577_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4576 N_OUT9_Mn9@4576_d N_OUT8_Mn9@4576_g N_VSS_Mn9@4576_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4577 N_OUT9_Mp9@4577_d N_OUT8_Mp9@4577_g N_VDD_Mp9@4577_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4576 N_OUT9_Mp9@4576_d N_OUT8_Mp9@4576_g N_VDD_Mp9@4576_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4575 N_OUT9_Mn9@4575_d N_OUT8_Mn9@4575_g N_VSS_Mn9@4575_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4574 N_OUT9_Mn9@4574_d N_OUT8_Mn9@4574_g N_VSS_Mn9@4574_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4575 N_OUT9_Mp9@4575_d N_OUT8_Mp9@4575_g N_VDD_Mp9@4575_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4574 N_OUT9_Mp9@4574_d N_OUT8_Mp9@4574_g N_VDD_Mp9@4574_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4573 N_OUT9_Mn9@4573_d N_OUT8_Mn9@4573_g N_VSS_Mn9@4573_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4572 N_OUT9_Mn9@4572_d N_OUT8_Mn9@4572_g N_VSS_Mn9@4572_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4573 N_OUT9_Mp9@4573_d N_OUT8_Mp9@4573_g N_VDD_Mp9@4573_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4572 N_OUT9_Mp9@4572_d N_OUT8_Mp9@4572_g N_VDD_Mp9@4572_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4571 N_OUT9_Mn9@4571_d N_OUT8_Mn9@4571_g N_VSS_Mn9@4571_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4570 N_OUT9_Mn9@4570_d N_OUT8_Mn9@4570_g N_VSS_Mn9@4570_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4571 N_OUT9_Mp9@4571_d N_OUT8_Mp9@4571_g N_VDD_Mp9@4571_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4570 N_OUT9_Mp9@4570_d N_OUT8_Mp9@4570_g N_VDD_Mp9@4570_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4569 N_OUT9_Mn9@4569_d N_OUT8_Mn9@4569_g N_VSS_Mn9@4569_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4568 N_OUT9_Mn9@4568_d N_OUT8_Mn9@4568_g N_VSS_Mn9@4568_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4569 N_OUT9_Mp9@4569_d N_OUT8_Mp9@4569_g N_VDD_Mp9@4569_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4568 N_OUT9_Mp9@4568_d N_OUT8_Mp9@4568_g N_VDD_Mp9@4568_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4567 N_OUT9_Mn9@4567_d N_OUT8_Mn9@4567_g N_VSS_Mn9@4567_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4566 N_OUT9_Mn9@4566_d N_OUT8_Mn9@4566_g N_VSS_Mn9@4566_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4567 N_OUT9_Mp9@4567_d N_OUT8_Mp9@4567_g N_VDD_Mp9@4567_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4566 N_OUT9_Mp9@4566_d N_OUT8_Mp9@4566_g N_VDD_Mp9@4566_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4565 N_OUT9_Mn9@4565_d N_OUT8_Mn9@4565_g N_VSS_Mn9@4565_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4564 N_OUT9_Mn9@4564_d N_OUT8_Mn9@4564_g N_VSS_Mn9@4564_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4565 N_OUT9_Mp9@4565_d N_OUT8_Mp9@4565_g N_VDD_Mp9@4565_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4564 N_OUT9_Mp9@4564_d N_OUT8_Mp9@4564_g N_VDD_Mp9@4564_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4563 N_OUT9_Mn9@4563_d N_OUT8_Mn9@4563_g N_VSS_Mn9@4563_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4562 N_OUT9_Mn9@4562_d N_OUT8_Mn9@4562_g N_VSS_Mn9@4562_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4563 N_OUT9_Mp9@4563_d N_OUT8_Mp9@4563_g N_VDD_Mp9@4563_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4562 N_OUT9_Mp9@4562_d N_OUT8_Mp9@4562_g N_VDD_Mp9@4562_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4561 N_OUT9_Mn9@4561_d N_OUT8_Mn9@4561_g N_VSS_Mn9@4561_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4560 N_OUT9_Mn9@4560_d N_OUT8_Mn9@4560_g N_VSS_Mn9@4560_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4561 N_OUT9_Mp9@4561_d N_OUT8_Mp9@4561_g N_VDD_Mp9@4561_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4560 N_OUT9_Mp9@4560_d N_OUT8_Mp9@4560_g N_VDD_Mp9@4560_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4559 N_OUT9_Mn9@4559_d N_OUT8_Mn9@4559_g N_VSS_Mn9@4559_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4558 N_OUT9_Mn9@4558_d N_OUT8_Mn9@4558_g N_VSS_Mn9@4558_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4559 N_OUT9_Mp9@4559_d N_OUT8_Mp9@4559_g N_VDD_Mp9@4559_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4558 N_OUT9_Mp9@4558_d N_OUT8_Mp9@4558_g N_VDD_Mp9@4558_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4557 N_OUT9_Mn9@4557_d N_OUT8_Mn9@4557_g N_VSS_Mn9@4557_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4556 N_OUT9_Mn9@4556_d N_OUT8_Mn9@4556_g N_VSS_Mn9@4556_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4557 N_OUT9_Mp9@4557_d N_OUT8_Mp9@4557_g N_VDD_Mp9@4557_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4556 N_OUT9_Mp9@4556_d N_OUT8_Mp9@4556_g N_VDD_Mp9@4556_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4555 N_OUT9_Mn9@4555_d N_OUT8_Mn9@4555_g N_VSS_Mn9@4555_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4554 N_OUT9_Mn9@4554_d N_OUT8_Mn9@4554_g N_VSS_Mn9@4554_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4555 N_OUT9_Mp9@4555_d N_OUT8_Mp9@4555_g N_VDD_Mp9@4555_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4554 N_OUT9_Mp9@4554_d N_OUT8_Mp9@4554_g N_VDD_Mp9@4554_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4553 N_OUT9_Mn9@4553_d N_OUT8_Mn9@4553_g N_VSS_Mn9@4553_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4552 N_OUT9_Mn9@4552_d N_OUT8_Mn9@4552_g N_VSS_Mn9@4552_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4553 N_OUT9_Mp9@4553_d N_OUT8_Mp9@4553_g N_VDD_Mp9@4553_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4552 N_OUT9_Mp9@4552_d N_OUT8_Mp9@4552_g N_VDD_Mp9@4552_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4551 N_OUT9_Mn9@4551_d N_OUT8_Mn9@4551_g N_VSS_Mn9@4551_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4550 N_OUT9_Mn9@4550_d N_OUT8_Mn9@4550_g N_VSS_Mn9@4550_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4551 N_OUT9_Mp9@4551_d N_OUT8_Mp9@4551_g N_VDD_Mp9@4551_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4550 N_OUT9_Mp9@4550_d N_OUT8_Mp9@4550_g N_VDD_Mp9@4550_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4549 N_OUT9_Mn9@4549_d N_OUT8_Mn9@4549_g N_VSS_Mn9@4549_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4548 N_OUT9_Mn9@4548_d N_OUT8_Mn9@4548_g N_VSS_Mn9@4548_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4549 N_OUT9_Mp9@4549_d N_OUT8_Mp9@4549_g N_VDD_Mp9@4549_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4548 N_OUT9_Mp9@4548_d N_OUT8_Mp9@4548_g N_VDD_Mp9@4548_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4547 N_OUT9_Mn9@4547_d N_OUT8_Mn9@4547_g N_VSS_Mn9@4547_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4546 N_OUT9_Mn9@4546_d N_OUT8_Mn9@4546_g N_VSS_Mn9@4546_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4547 N_OUT9_Mp9@4547_d N_OUT8_Mp9@4547_g N_VDD_Mp9@4547_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4546 N_OUT9_Mp9@4546_d N_OUT8_Mp9@4546_g N_VDD_Mp9@4546_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4545 N_OUT9_Mn9@4545_d N_OUT8_Mn9@4545_g N_VSS_Mn9@4545_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4544 N_OUT9_Mn9@4544_d N_OUT8_Mn9@4544_g N_VSS_Mn9@4544_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4545 N_OUT9_Mp9@4545_d N_OUT8_Mp9@4545_g N_VDD_Mp9@4545_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4544 N_OUT9_Mp9@4544_d N_OUT8_Mp9@4544_g N_VDD_Mp9@4544_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4543 N_OUT9_Mn9@4543_d N_OUT8_Mn9@4543_g N_VSS_Mn9@4543_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4542 N_OUT9_Mn9@4542_d N_OUT8_Mn9@4542_g N_VSS_Mn9@4542_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4543 N_OUT9_Mp9@4543_d N_OUT8_Mp9@4543_g N_VDD_Mp9@4543_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4542 N_OUT9_Mp9@4542_d N_OUT8_Mp9@4542_g N_VDD_Mp9@4542_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4541 N_OUT9_Mn9@4541_d N_OUT8_Mn9@4541_g N_VSS_Mn9@4541_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4540 N_OUT9_Mn9@4540_d N_OUT8_Mn9@4540_g N_VSS_Mn9@4540_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4541 N_OUT9_Mp9@4541_d N_OUT8_Mp9@4541_g N_VDD_Mp9@4541_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4540 N_OUT9_Mp9@4540_d N_OUT8_Mp9@4540_g N_VDD_Mp9@4540_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4539 N_OUT9_Mn9@4539_d N_OUT8_Mn9@4539_g N_VSS_Mn9@4539_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4538 N_OUT9_Mn9@4538_d N_OUT8_Mn9@4538_g N_VSS_Mn9@4538_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4539 N_OUT9_Mp9@4539_d N_OUT8_Mp9@4539_g N_VDD_Mp9@4539_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4538 N_OUT9_Mp9@4538_d N_OUT8_Mp9@4538_g N_VDD_Mp9@4538_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4537 N_OUT9_Mn9@4537_d N_OUT8_Mn9@4537_g N_VSS_Mn9@4537_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4536 N_OUT9_Mn9@4536_d N_OUT8_Mn9@4536_g N_VSS_Mn9@4536_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4537 N_OUT9_Mp9@4537_d N_OUT8_Mp9@4537_g N_VDD_Mp9@4537_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4536 N_OUT9_Mp9@4536_d N_OUT8_Mp9@4536_g N_VDD_Mp9@4536_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4535 N_OUT9_Mn9@4535_d N_OUT8_Mn9@4535_g N_VSS_Mn9@4535_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4534 N_OUT9_Mn9@4534_d N_OUT8_Mn9@4534_g N_VSS_Mn9@4534_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4535 N_OUT9_Mp9@4535_d N_OUT8_Mp9@4535_g N_VDD_Mp9@4535_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4534 N_OUT9_Mp9@4534_d N_OUT8_Mp9@4534_g N_VDD_Mp9@4534_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4533 N_OUT9_Mn9@4533_d N_OUT8_Mn9@4533_g N_VSS_Mn9@4533_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4532 N_OUT9_Mn9@4532_d N_OUT8_Mn9@4532_g N_VSS_Mn9@4532_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4533 N_OUT9_Mp9@4533_d N_OUT8_Mp9@4533_g N_VDD_Mp9@4533_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4532 N_OUT9_Mp9@4532_d N_OUT8_Mp9@4532_g N_VDD_Mp9@4532_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4531 N_OUT9_Mn9@4531_d N_OUT8_Mn9@4531_g N_VSS_Mn9@4531_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4530 N_OUT9_Mn9@4530_d N_OUT8_Mn9@4530_g N_VSS_Mn9@4530_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4531 N_OUT9_Mp9@4531_d N_OUT8_Mp9@4531_g N_VDD_Mp9@4531_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4530 N_OUT9_Mp9@4530_d N_OUT8_Mp9@4530_g N_VDD_Mp9@4530_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4529 N_OUT9_Mn9@4529_d N_OUT8_Mn9@4529_g N_VSS_Mn9@4529_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4528 N_OUT9_Mn9@4528_d N_OUT8_Mn9@4528_g N_VSS_Mn9@4528_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4529 N_OUT9_Mp9@4529_d N_OUT8_Mp9@4529_g N_VDD_Mp9@4529_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4528 N_OUT9_Mp9@4528_d N_OUT8_Mp9@4528_g N_VDD_Mp9@4528_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4527 N_OUT9_Mn9@4527_d N_OUT8_Mn9@4527_g N_VSS_Mn9@4527_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4526 N_OUT9_Mn9@4526_d N_OUT8_Mn9@4526_g N_VSS_Mn9@4526_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4527 N_OUT9_Mp9@4527_d N_OUT8_Mp9@4527_g N_VDD_Mp9@4527_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4526 N_OUT9_Mp9@4526_d N_OUT8_Mp9@4526_g N_VDD_Mp9@4526_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4525 N_OUT9_Mn9@4525_d N_OUT8_Mn9@4525_g N_VSS_Mn9@4525_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4524 N_OUT9_Mn9@4524_d N_OUT8_Mn9@4524_g N_VSS_Mn9@4524_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4525 N_OUT9_Mp9@4525_d N_OUT8_Mp9@4525_g N_VDD_Mp9@4525_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4524 N_OUT9_Mp9@4524_d N_OUT8_Mp9@4524_g N_VDD_Mp9@4524_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4523 N_OUT9_Mn9@4523_d N_OUT8_Mn9@4523_g N_VSS_Mn9@4523_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4522 N_OUT9_Mn9@4522_d N_OUT8_Mn9@4522_g N_VSS_Mn9@4522_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4523 N_OUT9_Mp9@4523_d N_OUT8_Mp9@4523_g N_VDD_Mp9@4523_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4522 N_OUT9_Mp9@4522_d N_OUT8_Mp9@4522_g N_VDD_Mp9@4522_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4521 N_OUT9_Mn9@4521_d N_OUT8_Mn9@4521_g N_VSS_Mn9@4521_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4520 N_OUT9_Mn9@4520_d N_OUT8_Mn9@4520_g N_VSS_Mn9@4520_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4521 N_OUT9_Mp9@4521_d N_OUT8_Mp9@4521_g N_VDD_Mp9@4521_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4520 N_OUT9_Mp9@4520_d N_OUT8_Mp9@4520_g N_VDD_Mp9@4520_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4519 N_OUT9_Mn9@4519_d N_OUT8_Mn9@4519_g N_VSS_Mn9@4519_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4518 N_OUT9_Mn9@4518_d N_OUT8_Mn9@4518_g N_VSS_Mn9@4518_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4519 N_OUT9_Mp9@4519_d N_OUT8_Mp9@4519_g N_VDD_Mp9@4519_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4518 N_OUT9_Mp9@4518_d N_OUT8_Mp9@4518_g N_VDD_Mp9@4518_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4517 N_OUT9_Mn9@4517_d N_OUT8_Mn9@4517_g N_VSS_Mn9@4517_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4516 N_OUT9_Mn9@4516_d N_OUT8_Mn9@4516_g N_VSS_Mn9@4516_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4517 N_OUT9_Mp9@4517_d N_OUT8_Mp9@4517_g N_VDD_Mp9@4517_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4516 N_OUT9_Mp9@4516_d N_OUT8_Mp9@4516_g N_VDD_Mp9@4516_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4515 N_OUT9_Mn9@4515_d N_OUT8_Mn9@4515_g N_VSS_Mn9@4515_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4514 N_OUT9_Mn9@4514_d N_OUT8_Mn9@4514_g N_VSS_Mn9@4514_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4515 N_OUT9_Mp9@4515_d N_OUT8_Mp9@4515_g N_VDD_Mp9@4515_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4514 N_OUT9_Mp9@4514_d N_OUT8_Mp9@4514_g N_VDD_Mp9@4514_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4513 N_OUT9_Mn9@4513_d N_OUT8_Mn9@4513_g N_VSS_Mn9@4513_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4512 N_OUT9_Mn9@4512_d N_OUT8_Mn9@4512_g N_VSS_Mn9@4512_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4513 N_OUT9_Mp9@4513_d N_OUT8_Mp9@4513_g N_VDD_Mp9@4513_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4512 N_OUT9_Mp9@4512_d N_OUT8_Mp9@4512_g N_VDD_Mp9@4512_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4511 N_OUT9_Mn9@4511_d N_OUT8_Mn9@4511_g N_VSS_Mn9@4511_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4510 N_OUT9_Mn9@4510_d N_OUT8_Mn9@4510_g N_VSS_Mn9@4510_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4511 N_OUT9_Mp9@4511_d N_OUT8_Mp9@4511_g N_VDD_Mp9@4511_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4510 N_OUT9_Mp9@4510_d N_OUT8_Mp9@4510_g N_VDD_Mp9@4510_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4509 N_OUT9_Mn9@4509_d N_OUT8_Mn9@4509_g N_VSS_Mn9@4509_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4508 N_OUT9_Mn9@4508_d N_OUT8_Mn9@4508_g N_VSS_Mn9@4508_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4509 N_OUT9_Mp9@4509_d N_OUT8_Mp9@4509_g N_VDD_Mp9@4509_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4508 N_OUT9_Mp9@4508_d N_OUT8_Mp9@4508_g N_VDD_Mp9@4508_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4507 N_OUT9_Mn9@4507_d N_OUT8_Mn9@4507_g N_VSS_Mn9@4507_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4506 N_OUT9_Mn9@4506_d N_OUT8_Mn9@4506_g N_VSS_Mn9@4506_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4507 N_OUT9_Mp9@4507_d N_OUT8_Mp9@4507_g N_VDD_Mp9@4507_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4506 N_OUT9_Mp9@4506_d N_OUT8_Mp9@4506_g N_VDD_Mp9@4506_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4505 N_OUT9_Mn9@4505_d N_OUT8_Mn9@4505_g N_VSS_Mn9@4505_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4504 N_OUT9_Mn9@4504_d N_OUT8_Mn9@4504_g N_VSS_Mn9@4504_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4505 N_OUT9_Mp9@4505_d N_OUT8_Mp9@4505_g N_VDD_Mp9@4505_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4504 N_OUT9_Mp9@4504_d N_OUT8_Mp9@4504_g N_VDD_Mp9@4504_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4503 N_OUT9_Mn9@4503_d N_OUT8_Mn9@4503_g N_VSS_Mn9@4503_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4502 N_OUT9_Mn9@4502_d N_OUT8_Mn9@4502_g N_VSS_Mn9@4502_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4503 N_OUT9_Mp9@4503_d N_OUT8_Mp9@4503_g N_VDD_Mp9@4503_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4502 N_OUT9_Mp9@4502_d N_OUT8_Mp9@4502_g N_VDD_Mp9@4502_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4501 N_OUT9_Mn9@4501_d N_OUT8_Mn9@4501_g N_VSS_Mn9@4501_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4500 N_OUT9_Mn9@4500_d N_OUT8_Mn9@4500_g N_VSS_Mn9@4500_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4501 N_OUT9_Mp9@4501_d N_OUT8_Mp9@4501_g N_VDD_Mp9@4501_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4500 N_OUT9_Mp9@4500_d N_OUT8_Mp9@4500_g N_VDD_Mp9@4500_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4499 N_OUT9_Mn9@4499_d N_OUT8_Mn9@4499_g N_VSS_Mn9@4499_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4498 N_OUT9_Mn9@4498_d N_OUT8_Mn9@4498_g N_VSS_Mn9@4498_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4499 N_OUT9_Mp9@4499_d N_OUT8_Mp9@4499_g N_VDD_Mp9@4499_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4498 N_OUT9_Mp9@4498_d N_OUT8_Mp9@4498_g N_VDD_Mp9@4498_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4497 N_OUT9_Mn9@4497_d N_OUT8_Mn9@4497_g N_VSS_Mn9@4497_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4496 N_OUT9_Mn9@4496_d N_OUT8_Mn9@4496_g N_VSS_Mn9@4496_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4497 N_OUT9_Mp9@4497_d N_OUT8_Mp9@4497_g N_VDD_Mp9@4497_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4496 N_OUT9_Mp9@4496_d N_OUT8_Mp9@4496_g N_VDD_Mp9@4496_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4495 N_OUT9_Mn9@4495_d N_OUT8_Mn9@4495_g N_VSS_Mn9@4495_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4494 N_OUT9_Mn9@4494_d N_OUT8_Mn9@4494_g N_VSS_Mn9@4494_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4495 N_OUT9_Mp9@4495_d N_OUT8_Mp9@4495_g N_VDD_Mp9@4495_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4494 N_OUT9_Mp9@4494_d N_OUT8_Mp9@4494_g N_VDD_Mp9@4494_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4493 N_OUT9_Mn9@4493_d N_OUT8_Mn9@4493_g N_VSS_Mn9@4493_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4492 N_OUT9_Mn9@4492_d N_OUT8_Mn9@4492_g N_VSS_Mn9@4492_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4493 N_OUT9_Mp9@4493_d N_OUT8_Mp9@4493_g N_VDD_Mp9@4493_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4492 N_OUT9_Mp9@4492_d N_OUT8_Mp9@4492_g N_VDD_Mp9@4492_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4491 N_OUT9_Mn9@4491_d N_OUT8_Mn9@4491_g N_VSS_Mn9@4491_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4490 N_OUT9_Mn9@4490_d N_OUT8_Mn9@4490_g N_VSS_Mn9@4490_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4491 N_OUT9_Mp9@4491_d N_OUT8_Mp9@4491_g N_VDD_Mp9@4491_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4490 N_OUT9_Mp9@4490_d N_OUT8_Mp9@4490_g N_VDD_Mp9@4490_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4489 N_OUT9_Mn9@4489_d N_OUT8_Mn9@4489_g N_VSS_Mn9@4489_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4488 N_OUT9_Mn9@4488_d N_OUT8_Mn9@4488_g N_VSS_Mn9@4488_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4489 N_OUT9_Mp9@4489_d N_OUT8_Mp9@4489_g N_VDD_Mp9@4489_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4488 N_OUT9_Mp9@4488_d N_OUT8_Mp9@4488_g N_VDD_Mp9@4488_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4487 N_OUT9_Mn9@4487_d N_OUT8_Mn9@4487_g N_VSS_Mn9@4487_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4486 N_OUT9_Mn9@4486_d N_OUT8_Mn9@4486_g N_VSS_Mn9@4486_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4487 N_OUT9_Mp9@4487_d N_OUT8_Mp9@4487_g N_VDD_Mp9@4487_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4486 N_OUT9_Mp9@4486_d N_OUT8_Mp9@4486_g N_VDD_Mp9@4486_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4485 N_OUT9_Mn9@4485_d N_OUT8_Mn9@4485_g N_VSS_Mn9@4485_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4484 N_OUT9_Mn9@4484_d N_OUT8_Mn9@4484_g N_VSS_Mn9@4484_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4485 N_OUT9_Mp9@4485_d N_OUT8_Mp9@4485_g N_VDD_Mp9@4485_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4484 N_OUT9_Mp9@4484_d N_OUT8_Mp9@4484_g N_VDD_Mp9@4484_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4483 N_OUT9_Mn9@4483_d N_OUT8_Mn9@4483_g N_VSS_Mn9@4483_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4482 N_OUT9_Mn9@4482_d N_OUT8_Mn9@4482_g N_VSS_Mn9@4482_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4483 N_OUT9_Mp9@4483_d N_OUT8_Mp9@4483_g N_VDD_Mp9@4483_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4482 N_OUT9_Mp9@4482_d N_OUT8_Mp9@4482_g N_VDD_Mp9@4482_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4481 N_OUT9_Mn9@4481_d N_OUT8_Mn9@4481_g N_VSS_Mn9@4481_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4480 N_OUT9_Mn9@4480_d N_OUT8_Mn9@4480_g N_VSS_Mn9@4480_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4481 N_OUT9_Mp9@4481_d N_OUT8_Mp9@4481_g N_VDD_Mp9@4481_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4480 N_OUT9_Mp9@4480_d N_OUT8_Mp9@4480_g N_VDD_Mp9@4480_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4479 N_OUT9_Mn9@4479_d N_OUT8_Mn9@4479_g N_VSS_Mn9@4479_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4478 N_OUT9_Mn9@4478_d N_OUT8_Mn9@4478_g N_VSS_Mn9@4478_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4479 N_OUT9_Mp9@4479_d N_OUT8_Mp9@4479_g N_VDD_Mp9@4479_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4478 N_OUT9_Mp9@4478_d N_OUT8_Mp9@4478_g N_VDD_Mp9@4478_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4477 N_OUT9_Mn9@4477_d N_OUT8_Mn9@4477_g N_VSS_Mn9@4477_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4476 N_OUT9_Mn9@4476_d N_OUT8_Mn9@4476_g N_VSS_Mn9@4476_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4477 N_OUT9_Mp9@4477_d N_OUT8_Mp9@4477_g N_VDD_Mp9@4477_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4476 N_OUT9_Mp9@4476_d N_OUT8_Mp9@4476_g N_VDD_Mp9@4476_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4475 N_OUT9_Mn9@4475_d N_OUT8_Mn9@4475_g N_VSS_Mn9@4475_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4474 N_OUT9_Mn9@4474_d N_OUT8_Mn9@4474_g N_VSS_Mn9@4474_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4475 N_OUT9_Mp9@4475_d N_OUT8_Mp9@4475_g N_VDD_Mp9@4475_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4474 N_OUT9_Mp9@4474_d N_OUT8_Mp9@4474_g N_VDD_Mp9@4474_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4473 N_OUT9_Mn9@4473_d N_OUT8_Mn9@4473_g N_VSS_Mn9@4473_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4472 N_OUT9_Mn9@4472_d N_OUT8_Mn9@4472_g N_VSS_Mn9@4472_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4473 N_OUT9_Mp9@4473_d N_OUT8_Mp9@4473_g N_VDD_Mp9@4473_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4472 N_OUT9_Mp9@4472_d N_OUT8_Mp9@4472_g N_VDD_Mp9@4472_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4471 N_OUT9_Mn9@4471_d N_OUT8_Mn9@4471_g N_VSS_Mn9@4471_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4470 N_OUT9_Mn9@4470_d N_OUT8_Mn9@4470_g N_VSS_Mn9@4470_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4471 N_OUT9_Mp9@4471_d N_OUT8_Mp9@4471_g N_VDD_Mp9@4471_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4470 N_OUT9_Mp9@4470_d N_OUT8_Mp9@4470_g N_VDD_Mp9@4470_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4469 N_OUT9_Mn9@4469_d N_OUT8_Mn9@4469_g N_VSS_Mn9@4469_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4468 N_OUT9_Mn9@4468_d N_OUT8_Mn9@4468_g N_VSS_Mn9@4468_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4469 N_OUT9_Mp9@4469_d N_OUT8_Mp9@4469_g N_VDD_Mp9@4469_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4468 N_OUT9_Mp9@4468_d N_OUT8_Mp9@4468_g N_VDD_Mp9@4468_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4467 N_OUT9_Mn9@4467_d N_OUT8_Mn9@4467_g N_VSS_Mn9@4467_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4466 N_OUT9_Mn9@4466_d N_OUT8_Mn9@4466_g N_VSS_Mn9@4466_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4467 N_OUT9_Mp9@4467_d N_OUT8_Mp9@4467_g N_VDD_Mp9@4467_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4466 N_OUT9_Mp9@4466_d N_OUT8_Mp9@4466_g N_VDD_Mp9@4466_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4465 N_OUT9_Mn9@4465_d N_OUT8_Mn9@4465_g N_VSS_Mn9@4465_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4464 N_OUT9_Mn9@4464_d N_OUT8_Mn9@4464_g N_VSS_Mn9@4464_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4465 N_OUT9_Mp9@4465_d N_OUT8_Mp9@4465_g N_VDD_Mp9@4465_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4464 N_OUT9_Mp9@4464_d N_OUT8_Mp9@4464_g N_VDD_Mp9@4464_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4463 N_OUT9_Mn9@4463_d N_OUT8_Mn9@4463_g N_VSS_Mn9@4463_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4462 N_OUT9_Mn9@4462_d N_OUT8_Mn9@4462_g N_VSS_Mn9@4462_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4463 N_OUT9_Mp9@4463_d N_OUT8_Mp9@4463_g N_VDD_Mp9@4463_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4462 N_OUT9_Mp9@4462_d N_OUT8_Mp9@4462_g N_VDD_Mp9@4462_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4461 N_OUT9_Mn9@4461_d N_OUT8_Mn9@4461_g N_VSS_Mn9@4461_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4460 N_OUT9_Mn9@4460_d N_OUT8_Mn9@4460_g N_VSS_Mn9@4460_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4461 N_OUT9_Mp9@4461_d N_OUT8_Mp9@4461_g N_VDD_Mp9@4461_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4460 N_OUT9_Mp9@4460_d N_OUT8_Mp9@4460_g N_VDD_Mp9@4460_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4459 N_OUT9_Mn9@4459_d N_OUT8_Mn9@4459_g N_VSS_Mn9@4459_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4458 N_OUT9_Mn9@4458_d N_OUT8_Mn9@4458_g N_VSS_Mn9@4458_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4459 N_OUT9_Mp9@4459_d N_OUT8_Mp9@4459_g N_VDD_Mp9@4459_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4458 N_OUT9_Mp9@4458_d N_OUT8_Mp9@4458_g N_VDD_Mp9@4458_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4457 N_OUT9_Mn9@4457_d N_OUT8_Mn9@4457_g N_VSS_Mn9@4457_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4456 N_OUT9_Mn9@4456_d N_OUT8_Mn9@4456_g N_VSS_Mn9@4456_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4457 N_OUT9_Mp9@4457_d N_OUT8_Mp9@4457_g N_VDD_Mp9@4457_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4456 N_OUT9_Mp9@4456_d N_OUT8_Mp9@4456_g N_VDD_Mp9@4456_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4455 N_OUT9_Mn9@4455_d N_OUT8_Mn9@4455_g N_VSS_Mn9@4455_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4454 N_OUT9_Mn9@4454_d N_OUT8_Mn9@4454_g N_VSS_Mn9@4454_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4455 N_OUT9_Mp9@4455_d N_OUT8_Mp9@4455_g N_VDD_Mp9@4455_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4454 N_OUT9_Mp9@4454_d N_OUT8_Mp9@4454_g N_VDD_Mp9@4454_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4453 N_OUT9_Mn9@4453_d N_OUT8_Mn9@4453_g N_VSS_Mn9@4453_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4452 N_OUT9_Mn9@4452_d N_OUT8_Mn9@4452_g N_VSS_Mn9@4452_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4453 N_OUT9_Mp9@4453_d N_OUT8_Mp9@4453_g N_VDD_Mp9@4453_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4452 N_OUT9_Mp9@4452_d N_OUT8_Mp9@4452_g N_VDD_Mp9@4452_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4451 N_OUT9_Mn9@4451_d N_OUT8_Mn9@4451_g N_VSS_Mn9@4451_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4450 N_OUT9_Mn9@4450_d N_OUT8_Mn9@4450_g N_VSS_Mn9@4450_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4451 N_OUT9_Mp9@4451_d N_OUT8_Mp9@4451_g N_VDD_Mp9@4451_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4450 N_OUT9_Mp9@4450_d N_OUT8_Mp9@4450_g N_VDD_Mp9@4450_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4449 N_OUT9_Mn9@4449_d N_OUT8_Mn9@4449_g N_VSS_Mn9@4449_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4448 N_OUT9_Mn9@4448_d N_OUT8_Mn9@4448_g N_VSS_Mn9@4448_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4449 N_OUT9_Mp9@4449_d N_OUT8_Mp9@4449_g N_VDD_Mp9@4449_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4448 N_OUT9_Mp9@4448_d N_OUT8_Mp9@4448_g N_VDD_Mp9@4448_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4447 N_OUT9_Mn9@4447_d N_OUT8_Mn9@4447_g N_VSS_Mn9@4447_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4446 N_OUT9_Mn9@4446_d N_OUT8_Mn9@4446_g N_VSS_Mn9@4446_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4447 N_OUT9_Mp9@4447_d N_OUT8_Mp9@4447_g N_VDD_Mp9@4447_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4446 N_OUT9_Mp9@4446_d N_OUT8_Mp9@4446_g N_VDD_Mp9@4446_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4445 N_OUT9_Mn9@4445_d N_OUT8_Mn9@4445_g N_VSS_Mn9@4445_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4444 N_OUT9_Mn9@4444_d N_OUT8_Mn9@4444_g N_VSS_Mn9@4444_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4445 N_OUT9_Mp9@4445_d N_OUT8_Mp9@4445_g N_VDD_Mp9@4445_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4444 N_OUT9_Mp9@4444_d N_OUT8_Mp9@4444_g N_VDD_Mp9@4444_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4443 N_OUT9_Mn9@4443_d N_OUT8_Mn9@4443_g N_VSS_Mn9@4443_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4442 N_OUT9_Mn9@4442_d N_OUT8_Mn9@4442_g N_VSS_Mn9@4442_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4443 N_OUT9_Mp9@4443_d N_OUT8_Mp9@4443_g N_VDD_Mp9@4443_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4442 N_OUT9_Mp9@4442_d N_OUT8_Mp9@4442_g N_VDD_Mp9@4442_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4441 N_OUT9_Mn9@4441_d N_OUT8_Mn9@4441_g N_VSS_Mn9@4441_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4440 N_OUT9_Mn9@4440_d N_OUT8_Mn9@4440_g N_VSS_Mn9@4440_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4441 N_OUT9_Mp9@4441_d N_OUT8_Mp9@4441_g N_VDD_Mp9@4441_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4440 N_OUT9_Mp9@4440_d N_OUT8_Mp9@4440_g N_VDD_Mp9@4440_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4439 N_OUT9_Mn9@4439_d N_OUT8_Mn9@4439_g N_VSS_Mn9@4439_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4438 N_OUT9_Mn9@4438_d N_OUT8_Mn9@4438_g N_VSS_Mn9@4438_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4439 N_OUT9_Mp9@4439_d N_OUT8_Mp9@4439_g N_VDD_Mp9@4439_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4438 N_OUT9_Mp9@4438_d N_OUT8_Mp9@4438_g N_VDD_Mp9@4438_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4437 N_OUT9_Mn9@4437_d N_OUT8_Mn9@4437_g N_VSS_Mn9@4437_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4436 N_OUT9_Mn9@4436_d N_OUT8_Mn9@4436_g N_VSS_Mn9@4436_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4437 N_OUT9_Mp9@4437_d N_OUT8_Mp9@4437_g N_VDD_Mp9@4437_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4436 N_OUT9_Mp9@4436_d N_OUT8_Mp9@4436_g N_VDD_Mp9@4436_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4435 N_OUT9_Mn9@4435_d N_OUT8_Mn9@4435_g N_VSS_Mn9@4435_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4434 N_OUT9_Mn9@4434_d N_OUT8_Mn9@4434_g N_VSS_Mn9@4434_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4435 N_OUT9_Mp9@4435_d N_OUT8_Mp9@4435_g N_VDD_Mp9@4435_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4434 N_OUT9_Mp9@4434_d N_OUT8_Mp9@4434_g N_VDD_Mp9@4434_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4433 N_OUT9_Mn9@4433_d N_OUT8_Mn9@4433_g N_VSS_Mn9@4433_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4432 N_OUT9_Mn9@4432_d N_OUT8_Mn9@4432_g N_VSS_Mn9@4432_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4433 N_OUT9_Mp9@4433_d N_OUT8_Mp9@4433_g N_VDD_Mp9@4433_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4432 N_OUT9_Mp9@4432_d N_OUT8_Mp9@4432_g N_VDD_Mp9@4432_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4431 N_OUT9_Mn9@4431_d N_OUT8_Mn9@4431_g N_VSS_Mn9@4431_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4430 N_OUT9_Mn9@4430_d N_OUT8_Mn9@4430_g N_VSS_Mn9@4430_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4431 N_OUT9_Mp9@4431_d N_OUT8_Mp9@4431_g N_VDD_Mp9@4431_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4430 N_OUT9_Mp9@4430_d N_OUT8_Mp9@4430_g N_VDD_Mp9@4430_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4429 N_OUT9_Mn9@4429_d N_OUT8_Mn9@4429_g N_VSS_Mn9@4429_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4428 N_OUT9_Mn9@4428_d N_OUT8_Mn9@4428_g N_VSS_Mn9@4428_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4429 N_OUT9_Mp9@4429_d N_OUT8_Mp9@4429_g N_VDD_Mp9@4429_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4428 N_OUT9_Mp9@4428_d N_OUT8_Mp9@4428_g N_VDD_Mp9@4428_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4427 N_OUT9_Mn9@4427_d N_OUT8_Mn9@4427_g N_VSS_Mn9@4427_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4426 N_OUT9_Mn9@4426_d N_OUT8_Mn9@4426_g N_VSS_Mn9@4426_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4427 N_OUT9_Mp9@4427_d N_OUT8_Mp9@4427_g N_VDD_Mp9@4427_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4426 N_OUT9_Mp9@4426_d N_OUT8_Mp9@4426_g N_VDD_Mp9@4426_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4425 N_OUT9_Mn9@4425_d N_OUT8_Mn9@4425_g N_VSS_Mn9@4425_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4424 N_OUT9_Mn9@4424_d N_OUT8_Mn9@4424_g N_VSS_Mn9@4424_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4425 N_OUT9_Mp9@4425_d N_OUT8_Mp9@4425_g N_VDD_Mp9@4425_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4424 N_OUT9_Mp9@4424_d N_OUT8_Mp9@4424_g N_VDD_Mp9@4424_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4423 N_OUT9_Mn9@4423_d N_OUT8_Mn9@4423_g N_VSS_Mn9@4423_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4422 N_OUT9_Mn9@4422_d N_OUT8_Mn9@4422_g N_VSS_Mn9@4422_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4423 N_OUT9_Mp9@4423_d N_OUT8_Mp9@4423_g N_VDD_Mp9@4423_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4422 N_OUT9_Mp9@4422_d N_OUT8_Mp9@4422_g N_VDD_Mp9@4422_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4421 N_OUT9_Mn9@4421_d N_OUT8_Mn9@4421_g N_VSS_Mn9@4421_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4420 N_OUT9_Mn9@4420_d N_OUT8_Mn9@4420_g N_VSS_Mn9@4420_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4421 N_OUT9_Mp9@4421_d N_OUT8_Mp9@4421_g N_VDD_Mp9@4421_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4420 N_OUT9_Mp9@4420_d N_OUT8_Mp9@4420_g N_VDD_Mp9@4420_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4419 N_OUT9_Mn9@4419_d N_OUT8_Mn9@4419_g N_VSS_Mn9@4419_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4418 N_OUT9_Mn9@4418_d N_OUT8_Mn9@4418_g N_VSS_Mn9@4418_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4419 N_OUT9_Mp9@4419_d N_OUT8_Mp9@4419_g N_VDD_Mp9@4419_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4418 N_OUT9_Mp9@4418_d N_OUT8_Mp9@4418_g N_VDD_Mp9@4418_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4417 N_OUT9_Mn9@4417_d N_OUT8_Mn9@4417_g N_VSS_Mn9@4417_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4416 N_OUT9_Mn9@4416_d N_OUT8_Mn9@4416_g N_VSS_Mn9@4416_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4417 N_OUT9_Mp9@4417_d N_OUT8_Mp9@4417_g N_VDD_Mp9@4417_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4416 N_OUT9_Mp9@4416_d N_OUT8_Mp9@4416_g N_VDD_Mp9@4416_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4415 N_OUT9_Mn9@4415_d N_OUT8_Mn9@4415_g N_VSS_Mn9@4415_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4414 N_OUT9_Mn9@4414_d N_OUT8_Mn9@4414_g N_VSS_Mn9@4414_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4415 N_OUT9_Mp9@4415_d N_OUT8_Mp9@4415_g N_VDD_Mp9@4415_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4414 N_OUT9_Mp9@4414_d N_OUT8_Mp9@4414_g N_VDD_Mp9@4414_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4413 N_OUT9_Mn9@4413_d N_OUT8_Mn9@4413_g N_VSS_Mn9@4413_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4412 N_OUT9_Mn9@4412_d N_OUT8_Mn9@4412_g N_VSS_Mn9@4412_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4413 N_OUT9_Mp9@4413_d N_OUT8_Mp9@4413_g N_VDD_Mp9@4413_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4412 N_OUT9_Mp9@4412_d N_OUT8_Mp9@4412_g N_VDD_Mp9@4412_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4411 N_OUT9_Mn9@4411_d N_OUT8_Mn9@4411_g N_VSS_Mn9@4411_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4410 N_OUT9_Mn9@4410_d N_OUT8_Mn9@4410_g N_VSS_Mn9@4410_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4411 N_OUT9_Mp9@4411_d N_OUT8_Mp9@4411_g N_VDD_Mp9@4411_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4410 N_OUT9_Mp9@4410_d N_OUT8_Mp9@4410_g N_VDD_Mp9@4410_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4409 N_OUT9_Mn9@4409_d N_OUT8_Mn9@4409_g N_VSS_Mn9@4409_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4408 N_OUT9_Mn9@4408_d N_OUT8_Mn9@4408_g N_VSS_Mn9@4408_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4409 N_OUT9_Mp9@4409_d N_OUT8_Mp9@4409_g N_VDD_Mp9@4409_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4408 N_OUT9_Mp9@4408_d N_OUT8_Mp9@4408_g N_VDD_Mp9@4408_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4407 N_OUT9_Mn9@4407_d N_OUT8_Mn9@4407_g N_VSS_Mn9@4407_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4406 N_OUT9_Mn9@4406_d N_OUT8_Mn9@4406_g N_VSS_Mn9@4406_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4407 N_OUT9_Mp9@4407_d N_OUT8_Mp9@4407_g N_VDD_Mp9@4407_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4406 N_OUT9_Mp9@4406_d N_OUT8_Mp9@4406_g N_VDD_Mp9@4406_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4405 N_OUT9_Mn9@4405_d N_OUT8_Mn9@4405_g N_VSS_Mn9@4405_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4404 N_OUT9_Mn9@4404_d N_OUT8_Mn9@4404_g N_VSS_Mn9@4404_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4405 N_OUT9_Mp9@4405_d N_OUT8_Mp9@4405_g N_VDD_Mp9@4405_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4404 N_OUT9_Mp9@4404_d N_OUT8_Mp9@4404_g N_VDD_Mp9@4404_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4403 N_OUT9_Mn9@4403_d N_OUT8_Mn9@4403_g N_VSS_Mn9@4403_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4402 N_OUT9_Mn9@4402_d N_OUT8_Mn9@4402_g N_VSS_Mn9@4402_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4403 N_OUT9_Mp9@4403_d N_OUT8_Mp9@4403_g N_VDD_Mp9@4403_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4402 N_OUT9_Mp9@4402_d N_OUT8_Mp9@4402_g N_VDD_Mp9@4402_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4401 N_OUT9_Mn9@4401_d N_OUT8_Mn9@4401_g N_VSS_Mn9@4401_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4400 N_OUT9_Mn9@4400_d N_OUT8_Mn9@4400_g N_VSS_Mn9@4400_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4401 N_OUT9_Mp9@4401_d N_OUT8_Mp9@4401_g N_VDD_Mp9@4401_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4400 N_OUT9_Mp9@4400_d N_OUT8_Mp9@4400_g N_VDD_Mp9@4400_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4399 N_OUT9_Mn9@4399_d N_OUT8_Mn9@4399_g N_VSS_Mn9@4399_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4398 N_OUT9_Mn9@4398_d N_OUT8_Mn9@4398_g N_VSS_Mn9@4398_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4399 N_OUT9_Mp9@4399_d N_OUT8_Mp9@4399_g N_VDD_Mp9@4399_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4398 N_OUT9_Mp9@4398_d N_OUT8_Mp9@4398_g N_VDD_Mp9@4398_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4397 N_OUT9_Mn9@4397_d N_OUT8_Mn9@4397_g N_VSS_Mn9@4397_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4396 N_OUT9_Mn9@4396_d N_OUT8_Mn9@4396_g N_VSS_Mn9@4396_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4397 N_OUT9_Mp9@4397_d N_OUT8_Mp9@4397_g N_VDD_Mp9@4397_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4396 N_OUT9_Mp9@4396_d N_OUT8_Mp9@4396_g N_VDD_Mp9@4396_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4395 N_OUT9_Mn9@4395_d N_OUT8_Mn9@4395_g N_VSS_Mn9@4395_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4394 N_OUT9_Mn9@4394_d N_OUT8_Mn9@4394_g N_VSS_Mn9@4394_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4395 N_OUT9_Mp9@4395_d N_OUT8_Mp9@4395_g N_VDD_Mp9@4395_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4394 N_OUT9_Mp9@4394_d N_OUT8_Mp9@4394_g N_VDD_Mp9@4394_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4393 N_OUT9_Mn9@4393_d N_OUT8_Mn9@4393_g N_VSS_Mn9@4393_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4392 N_OUT9_Mn9@4392_d N_OUT8_Mn9@4392_g N_VSS_Mn9@4392_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4393 N_OUT9_Mp9@4393_d N_OUT8_Mp9@4393_g N_VDD_Mp9@4393_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4392 N_OUT9_Mp9@4392_d N_OUT8_Mp9@4392_g N_VDD_Mp9@4392_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4391 N_OUT9_Mn9@4391_d N_OUT8_Mn9@4391_g N_VSS_Mn9@4391_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4390 N_OUT9_Mn9@4390_d N_OUT8_Mn9@4390_g N_VSS_Mn9@4390_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4391 N_OUT9_Mp9@4391_d N_OUT8_Mp9@4391_g N_VDD_Mp9@4391_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4390 N_OUT9_Mp9@4390_d N_OUT8_Mp9@4390_g N_VDD_Mp9@4390_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4389 N_OUT9_Mn9@4389_d N_OUT8_Mn9@4389_g N_VSS_Mn9@4389_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4388 N_OUT9_Mn9@4388_d N_OUT8_Mn9@4388_g N_VSS_Mn9@4388_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4389 N_OUT9_Mp9@4389_d N_OUT8_Mp9@4389_g N_VDD_Mp9@4389_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4388 N_OUT9_Mp9@4388_d N_OUT8_Mp9@4388_g N_VDD_Mp9@4388_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4387 N_OUT9_Mn9@4387_d N_OUT8_Mn9@4387_g N_VSS_Mn9@4387_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4386 N_OUT9_Mn9@4386_d N_OUT8_Mn9@4386_g N_VSS_Mn9@4386_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4387 N_OUT9_Mp9@4387_d N_OUT8_Mp9@4387_g N_VDD_Mp9@4387_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4386 N_OUT9_Mp9@4386_d N_OUT8_Mp9@4386_g N_VDD_Mp9@4386_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4385 N_OUT9_Mn9@4385_d N_OUT8_Mn9@4385_g N_VSS_Mn9@4385_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4384 N_OUT9_Mn9@4384_d N_OUT8_Mn9@4384_g N_VSS_Mn9@4384_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4385 N_OUT9_Mp9@4385_d N_OUT8_Mp9@4385_g N_VDD_Mp9@4385_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4384 N_OUT9_Mp9@4384_d N_OUT8_Mp9@4384_g N_VDD_Mp9@4384_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4383 N_OUT9_Mn9@4383_d N_OUT8_Mn9@4383_g N_VSS_Mn9@4383_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4382 N_OUT9_Mn9@4382_d N_OUT8_Mn9@4382_g N_VSS_Mn9@4382_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4383 N_OUT9_Mp9@4383_d N_OUT8_Mp9@4383_g N_VDD_Mp9@4383_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4382 N_OUT9_Mp9@4382_d N_OUT8_Mp9@4382_g N_VDD_Mp9@4382_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4381 N_OUT9_Mn9@4381_d N_OUT8_Mn9@4381_g N_VSS_Mn9@4381_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4380 N_OUT9_Mn9@4380_d N_OUT8_Mn9@4380_g N_VSS_Mn9@4380_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4381 N_OUT9_Mp9@4381_d N_OUT8_Mp9@4381_g N_VDD_Mp9@4381_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4380 N_OUT9_Mp9@4380_d N_OUT8_Mp9@4380_g N_VDD_Mp9@4380_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4379 N_OUT9_Mn9@4379_d N_OUT8_Mn9@4379_g N_VSS_Mn9@4379_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4378 N_OUT9_Mn9@4378_d N_OUT8_Mn9@4378_g N_VSS_Mn9@4378_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4379 N_OUT9_Mp9@4379_d N_OUT8_Mp9@4379_g N_VDD_Mp9@4379_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4378 N_OUT9_Mp9@4378_d N_OUT8_Mp9@4378_g N_VDD_Mp9@4378_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4377 N_OUT9_Mn9@4377_d N_OUT8_Mn9@4377_g N_VSS_Mn9@4377_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4376 N_OUT9_Mn9@4376_d N_OUT8_Mn9@4376_g N_VSS_Mn9@4376_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4377 N_OUT9_Mp9@4377_d N_OUT8_Mp9@4377_g N_VDD_Mp9@4377_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4376 N_OUT9_Mp9@4376_d N_OUT8_Mp9@4376_g N_VDD_Mp9@4376_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4375 N_OUT9_Mn9@4375_d N_OUT8_Mn9@4375_g N_VSS_Mn9@4375_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4374 N_OUT9_Mn9@4374_d N_OUT8_Mn9@4374_g N_VSS_Mn9@4374_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4375 N_OUT9_Mp9@4375_d N_OUT8_Mp9@4375_g N_VDD_Mp9@4375_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4374 N_OUT9_Mp9@4374_d N_OUT8_Mp9@4374_g N_VDD_Mp9@4374_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4373 N_OUT9_Mn9@4373_d N_OUT8_Mn9@4373_g N_VSS_Mn9@4373_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4372 N_OUT9_Mn9@4372_d N_OUT8_Mn9@4372_g N_VSS_Mn9@4372_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4373 N_OUT9_Mp9@4373_d N_OUT8_Mp9@4373_g N_VDD_Mp9@4373_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4372 N_OUT9_Mp9@4372_d N_OUT8_Mp9@4372_g N_VDD_Mp9@4372_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4371 N_OUT9_Mn9@4371_d N_OUT8_Mn9@4371_g N_VSS_Mn9@4371_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4370 N_OUT9_Mn9@4370_d N_OUT8_Mn9@4370_g N_VSS_Mn9@4370_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4371 N_OUT9_Mp9@4371_d N_OUT8_Mp9@4371_g N_VDD_Mp9@4371_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4370 N_OUT9_Mp9@4370_d N_OUT8_Mp9@4370_g N_VDD_Mp9@4370_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4369 N_OUT9_Mn9@4369_d N_OUT8_Mn9@4369_g N_VSS_Mn9@4369_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4368 N_OUT9_Mn9@4368_d N_OUT8_Mn9@4368_g N_VSS_Mn9@4368_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4369 N_OUT9_Mp9@4369_d N_OUT8_Mp9@4369_g N_VDD_Mp9@4369_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4368 N_OUT9_Mp9@4368_d N_OUT8_Mp9@4368_g N_VDD_Mp9@4368_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4367 N_OUT9_Mn9@4367_d N_OUT8_Mn9@4367_g N_VSS_Mn9@4367_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4366 N_OUT9_Mn9@4366_d N_OUT8_Mn9@4366_g N_VSS_Mn9@4366_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4367 N_OUT9_Mp9@4367_d N_OUT8_Mp9@4367_g N_VDD_Mp9@4367_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4366 N_OUT9_Mp9@4366_d N_OUT8_Mp9@4366_g N_VDD_Mp9@4366_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4365 N_OUT9_Mn9@4365_d N_OUT8_Mn9@4365_g N_VSS_Mn9@4365_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4364 N_OUT9_Mn9@4364_d N_OUT8_Mn9@4364_g N_VSS_Mn9@4364_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4365 N_OUT9_Mp9@4365_d N_OUT8_Mp9@4365_g N_VDD_Mp9@4365_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4364 N_OUT9_Mp9@4364_d N_OUT8_Mp9@4364_g N_VDD_Mp9@4364_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4363 N_OUT9_Mn9@4363_d N_OUT8_Mn9@4363_g N_VSS_Mn9@4363_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4362 N_OUT9_Mn9@4362_d N_OUT8_Mn9@4362_g N_VSS_Mn9@4362_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4363 N_OUT9_Mp9@4363_d N_OUT8_Mp9@4363_g N_VDD_Mp9@4363_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4362 N_OUT9_Mp9@4362_d N_OUT8_Mp9@4362_g N_VDD_Mp9@4362_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4361 N_OUT9_Mn9@4361_d N_OUT8_Mn9@4361_g N_VSS_Mn9@4361_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4360 N_OUT9_Mn9@4360_d N_OUT8_Mn9@4360_g N_VSS_Mn9@4360_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4361 N_OUT9_Mp9@4361_d N_OUT8_Mp9@4361_g N_VDD_Mp9@4361_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4360 N_OUT9_Mp9@4360_d N_OUT8_Mp9@4360_g N_VDD_Mp9@4360_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4359 N_OUT9_Mn9@4359_d N_OUT8_Mn9@4359_g N_VSS_Mn9@4359_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4358 N_OUT9_Mn9@4358_d N_OUT8_Mn9@4358_g N_VSS_Mn9@4358_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4359 N_OUT9_Mp9@4359_d N_OUT8_Mp9@4359_g N_VDD_Mp9@4359_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4358 N_OUT9_Mp9@4358_d N_OUT8_Mp9@4358_g N_VDD_Mp9@4358_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4357 N_OUT9_Mn9@4357_d N_OUT8_Mn9@4357_g N_VSS_Mn9@4357_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4356 N_OUT9_Mn9@4356_d N_OUT8_Mn9@4356_g N_VSS_Mn9@4356_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4357 N_OUT9_Mp9@4357_d N_OUT8_Mp9@4357_g N_VDD_Mp9@4357_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4356 N_OUT9_Mp9@4356_d N_OUT8_Mp9@4356_g N_VDD_Mp9@4356_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4355 N_OUT9_Mn9@4355_d N_OUT8_Mn9@4355_g N_VSS_Mn9@4355_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4354 N_OUT9_Mn9@4354_d N_OUT8_Mn9@4354_g N_VSS_Mn9@4354_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4355 N_OUT9_Mp9@4355_d N_OUT8_Mp9@4355_g N_VDD_Mp9@4355_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4354 N_OUT9_Mp9@4354_d N_OUT8_Mp9@4354_g N_VDD_Mp9@4354_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4353 N_OUT9_Mn9@4353_d N_OUT8_Mn9@4353_g N_VSS_Mn9@4353_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4352 N_OUT9_Mn9@4352_d N_OUT8_Mn9@4352_g N_VSS_Mn9@4352_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4353 N_OUT9_Mp9@4353_d N_OUT8_Mp9@4353_g N_VDD_Mp9@4353_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4352 N_OUT9_Mp9@4352_d N_OUT8_Mp9@4352_g N_VDD_Mp9@4352_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4351 N_OUT9_Mn9@4351_d N_OUT8_Mn9@4351_g N_VSS_Mn9@4351_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4350 N_OUT9_Mn9@4350_d N_OUT8_Mn9@4350_g N_VSS_Mn9@4350_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4351 N_OUT9_Mp9@4351_d N_OUT8_Mp9@4351_g N_VDD_Mp9@4351_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4350 N_OUT9_Mp9@4350_d N_OUT8_Mp9@4350_g N_VDD_Mp9@4350_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4349 N_OUT9_Mn9@4349_d N_OUT8_Mn9@4349_g N_VSS_Mn9@4349_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4348 N_OUT9_Mn9@4348_d N_OUT8_Mn9@4348_g N_VSS_Mn9@4348_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4349 N_OUT9_Mp9@4349_d N_OUT8_Mp9@4349_g N_VDD_Mp9@4349_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4348 N_OUT9_Mp9@4348_d N_OUT8_Mp9@4348_g N_VDD_Mp9@4348_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4347 N_OUT9_Mn9@4347_d N_OUT8_Mn9@4347_g N_VSS_Mn9@4347_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4346 N_OUT9_Mn9@4346_d N_OUT8_Mn9@4346_g N_VSS_Mn9@4346_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4347 N_OUT9_Mp9@4347_d N_OUT8_Mp9@4347_g N_VDD_Mp9@4347_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4346 N_OUT9_Mp9@4346_d N_OUT8_Mp9@4346_g N_VDD_Mp9@4346_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4345 N_OUT9_Mn9@4345_d N_OUT8_Mn9@4345_g N_VSS_Mn9@4345_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4344 N_OUT9_Mn9@4344_d N_OUT8_Mn9@4344_g N_VSS_Mn9@4344_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4345 N_OUT9_Mp9@4345_d N_OUT8_Mp9@4345_g N_VDD_Mp9@4345_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4344 N_OUT9_Mp9@4344_d N_OUT8_Mp9@4344_g N_VDD_Mp9@4344_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4343 N_OUT9_Mn9@4343_d N_OUT8_Mn9@4343_g N_VSS_Mn9@4343_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4342 N_OUT9_Mn9@4342_d N_OUT8_Mn9@4342_g N_VSS_Mn9@4342_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4343 N_OUT9_Mp9@4343_d N_OUT8_Mp9@4343_g N_VDD_Mp9@4343_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4342 N_OUT9_Mp9@4342_d N_OUT8_Mp9@4342_g N_VDD_Mp9@4342_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4341 N_OUT9_Mn9@4341_d N_OUT8_Mn9@4341_g N_VSS_Mn9@4341_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4340 N_OUT9_Mn9@4340_d N_OUT8_Mn9@4340_g N_VSS_Mn9@4340_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4341 N_OUT9_Mp9@4341_d N_OUT8_Mp9@4341_g N_VDD_Mp9@4341_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4340 N_OUT9_Mp9@4340_d N_OUT8_Mp9@4340_g N_VDD_Mp9@4340_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4339 N_OUT9_Mn9@4339_d N_OUT8_Mn9@4339_g N_VSS_Mn9@4339_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4338 N_OUT9_Mn9@4338_d N_OUT8_Mn9@4338_g N_VSS_Mn9@4338_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4339 N_OUT9_Mp9@4339_d N_OUT8_Mp9@4339_g N_VDD_Mp9@4339_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4338 N_OUT9_Mp9@4338_d N_OUT8_Mp9@4338_g N_VDD_Mp9@4338_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4337 N_OUT9_Mn9@4337_d N_OUT8_Mn9@4337_g N_VSS_Mn9@4337_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4336 N_OUT9_Mn9@4336_d N_OUT8_Mn9@4336_g N_VSS_Mn9@4336_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4337 N_OUT9_Mp9@4337_d N_OUT8_Mp9@4337_g N_VDD_Mp9@4337_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4336 N_OUT9_Mp9@4336_d N_OUT8_Mp9@4336_g N_VDD_Mp9@4336_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4335 N_OUT9_Mn9@4335_d N_OUT8_Mn9@4335_g N_VSS_Mn9@4335_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4334 N_OUT9_Mn9@4334_d N_OUT8_Mn9@4334_g N_VSS_Mn9@4334_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4335 N_OUT9_Mp9@4335_d N_OUT8_Mp9@4335_g N_VDD_Mp9@4335_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4334 N_OUT9_Mp9@4334_d N_OUT8_Mp9@4334_g N_VDD_Mp9@4334_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4333 N_OUT9_Mn9@4333_d N_OUT8_Mn9@4333_g N_VSS_Mn9@4333_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4332 N_OUT9_Mn9@4332_d N_OUT8_Mn9@4332_g N_VSS_Mn9@4332_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4333 N_OUT9_Mp9@4333_d N_OUT8_Mp9@4333_g N_VDD_Mp9@4333_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4332 N_OUT9_Mp9@4332_d N_OUT8_Mp9@4332_g N_VDD_Mp9@4332_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4331 N_OUT9_Mn9@4331_d N_OUT8_Mn9@4331_g N_VSS_Mn9@4331_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4330 N_OUT9_Mn9@4330_d N_OUT8_Mn9@4330_g N_VSS_Mn9@4330_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4331 N_OUT9_Mp9@4331_d N_OUT8_Mp9@4331_g N_VDD_Mp9@4331_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4330 N_OUT9_Mp9@4330_d N_OUT8_Mp9@4330_g N_VDD_Mp9@4330_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4329 N_OUT9_Mn9@4329_d N_OUT8_Mn9@4329_g N_VSS_Mn9@4329_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4328 N_OUT9_Mn9@4328_d N_OUT8_Mn9@4328_g N_VSS_Mn9@4328_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4329 N_OUT9_Mp9@4329_d N_OUT8_Mp9@4329_g N_VDD_Mp9@4329_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4328 N_OUT9_Mp9@4328_d N_OUT8_Mp9@4328_g N_VDD_Mp9@4328_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4327 N_OUT9_Mn9@4327_d N_OUT8_Mn9@4327_g N_VSS_Mn9@4327_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4326 N_OUT9_Mn9@4326_d N_OUT8_Mn9@4326_g N_VSS_Mn9@4326_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4327 N_OUT9_Mp9@4327_d N_OUT8_Mp9@4327_g N_VDD_Mp9@4327_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4326 N_OUT9_Mp9@4326_d N_OUT8_Mp9@4326_g N_VDD_Mp9@4326_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4325 N_OUT9_Mn9@4325_d N_OUT8_Mn9@4325_g N_VSS_Mn9@4325_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4324 N_OUT9_Mn9@4324_d N_OUT8_Mn9@4324_g N_VSS_Mn9@4324_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4325 N_OUT9_Mp9@4325_d N_OUT8_Mp9@4325_g N_VDD_Mp9@4325_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4324 N_OUT9_Mp9@4324_d N_OUT8_Mp9@4324_g N_VDD_Mp9@4324_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4323 N_OUT9_Mn9@4323_d N_OUT8_Mn9@4323_g N_VSS_Mn9@4323_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4322 N_OUT9_Mn9@4322_d N_OUT8_Mn9@4322_g N_VSS_Mn9@4322_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4323 N_OUT9_Mp9@4323_d N_OUT8_Mp9@4323_g N_VDD_Mp9@4323_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4322 N_OUT9_Mp9@4322_d N_OUT8_Mp9@4322_g N_VDD_Mp9@4322_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4321 N_OUT9_Mn9@4321_d N_OUT8_Mn9@4321_g N_VSS_Mn9@4321_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4320 N_OUT9_Mn9@4320_d N_OUT8_Mn9@4320_g N_VSS_Mn9@4320_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4321 N_OUT9_Mp9@4321_d N_OUT8_Mp9@4321_g N_VDD_Mp9@4321_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4320 N_OUT9_Mp9@4320_d N_OUT8_Mp9@4320_g N_VDD_Mp9@4320_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4319 N_OUT9_Mn9@4319_d N_OUT8_Mn9@4319_g N_VSS_Mn9@4319_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4318 N_OUT9_Mn9@4318_d N_OUT8_Mn9@4318_g N_VSS_Mn9@4318_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4319 N_OUT9_Mp9@4319_d N_OUT8_Mp9@4319_g N_VDD_Mp9@4319_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4318 N_OUT9_Mp9@4318_d N_OUT8_Mp9@4318_g N_VDD_Mp9@4318_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4317 N_OUT9_Mn9@4317_d N_OUT8_Mn9@4317_g N_VSS_Mn9@4317_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4316 N_OUT9_Mn9@4316_d N_OUT8_Mn9@4316_g N_VSS_Mn9@4316_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4317 N_OUT9_Mp9@4317_d N_OUT8_Mp9@4317_g N_VDD_Mp9@4317_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4316 N_OUT9_Mp9@4316_d N_OUT8_Mp9@4316_g N_VDD_Mp9@4316_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4315 N_OUT9_Mn9@4315_d N_OUT8_Mn9@4315_g N_VSS_Mn9@4315_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4314 N_OUT9_Mn9@4314_d N_OUT8_Mn9@4314_g N_VSS_Mn9@4314_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4315 N_OUT9_Mp9@4315_d N_OUT8_Mp9@4315_g N_VDD_Mp9@4315_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4314 N_OUT9_Mp9@4314_d N_OUT8_Mp9@4314_g N_VDD_Mp9@4314_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4313 N_OUT9_Mn9@4313_d N_OUT8_Mn9@4313_g N_VSS_Mn9@4313_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4312 N_OUT9_Mn9@4312_d N_OUT8_Mn9@4312_g N_VSS_Mn9@4312_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4313 N_OUT9_Mp9@4313_d N_OUT8_Mp9@4313_g N_VDD_Mp9@4313_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4312 N_OUT9_Mp9@4312_d N_OUT8_Mp9@4312_g N_VDD_Mp9@4312_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4311 N_OUT9_Mn9@4311_d N_OUT8_Mn9@4311_g N_VSS_Mn9@4311_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4310 N_OUT9_Mn9@4310_d N_OUT8_Mn9@4310_g N_VSS_Mn9@4310_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4311 N_OUT9_Mp9@4311_d N_OUT8_Mp9@4311_g N_VDD_Mp9@4311_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4310 N_OUT9_Mp9@4310_d N_OUT8_Mp9@4310_g N_VDD_Mp9@4310_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4309 N_OUT9_Mn9@4309_d N_OUT8_Mn9@4309_g N_VSS_Mn9@4309_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4308 N_OUT9_Mn9@4308_d N_OUT8_Mn9@4308_g N_VSS_Mn9@4308_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4309 N_OUT9_Mp9@4309_d N_OUT8_Mp9@4309_g N_VDD_Mp9@4309_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4308 N_OUT9_Mp9@4308_d N_OUT8_Mp9@4308_g N_VDD_Mp9@4308_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4307 N_OUT9_Mn9@4307_d N_OUT8_Mn9@4307_g N_VSS_Mn9@4307_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4306 N_OUT9_Mn9@4306_d N_OUT8_Mn9@4306_g N_VSS_Mn9@4306_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4307 N_OUT9_Mp9@4307_d N_OUT8_Mp9@4307_g N_VDD_Mp9@4307_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4306 N_OUT9_Mp9@4306_d N_OUT8_Mp9@4306_g N_VDD_Mp9@4306_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4305 N_OUT9_Mn9@4305_d N_OUT8_Mn9@4305_g N_VSS_Mn9@4305_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4304 N_OUT9_Mn9@4304_d N_OUT8_Mn9@4304_g N_VSS_Mn9@4304_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4305 N_OUT9_Mp9@4305_d N_OUT8_Mp9@4305_g N_VDD_Mp9@4305_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4304 N_OUT9_Mp9@4304_d N_OUT8_Mp9@4304_g N_VDD_Mp9@4304_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4303 N_OUT9_Mn9@4303_d N_OUT8_Mn9@4303_g N_VSS_Mn9@4303_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4302 N_OUT9_Mn9@4302_d N_OUT8_Mn9@4302_g N_VSS_Mn9@4302_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4303 N_OUT9_Mp9@4303_d N_OUT8_Mp9@4303_g N_VDD_Mp9@4303_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4302 N_OUT9_Mp9@4302_d N_OUT8_Mp9@4302_g N_VDD_Mp9@4302_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4301 N_OUT9_Mn9@4301_d N_OUT8_Mn9@4301_g N_VSS_Mn9@4301_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4300 N_OUT9_Mn9@4300_d N_OUT8_Mn9@4300_g N_VSS_Mn9@4300_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4301 N_OUT9_Mp9@4301_d N_OUT8_Mp9@4301_g N_VDD_Mp9@4301_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4300 N_OUT9_Mp9@4300_d N_OUT8_Mp9@4300_g N_VDD_Mp9@4300_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4299 N_OUT9_Mn9@4299_d N_OUT8_Mn9@4299_g N_VSS_Mn9@4299_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4298 N_OUT9_Mn9@4298_d N_OUT8_Mn9@4298_g N_VSS_Mn9@4298_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4299 N_OUT9_Mp9@4299_d N_OUT8_Mp9@4299_g N_VDD_Mp9@4299_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4298 N_OUT9_Mp9@4298_d N_OUT8_Mp9@4298_g N_VDD_Mp9@4298_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4297 N_OUT9_Mn9@4297_d N_OUT8_Mn9@4297_g N_VSS_Mn9@4297_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4296 N_OUT9_Mn9@4296_d N_OUT8_Mn9@4296_g N_VSS_Mn9@4296_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4297 N_OUT9_Mp9@4297_d N_OUT8_Mp9@4297_g N_VDD_Mp9@4297_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4296 N_OUT9_Mp9@4296_d N_OUT8_Mp9@4296_g N_VDD_Mp9@4296_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4295 N_OUT9_Mn9@4295_d N_OUT8_Mn9@4295_g N_VSS_Mn9@4295_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4294 N_OUT9_Mn9@4294_d N_OUT8_Mn9@4294_g N_VSS_Mn9@4294_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4295 N_OUT9_Mp9@4295_d N_OUT8_Mp9@4295_g N_VDD_Mp9@4295_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4294 N_OUT9_Mp9@4294_d N_OUT8_Mp9@4294_g N_VDD_Mp9@4294_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4293 N_OUT9_Mn9@4293_d N_OUT8_Mn9@4293_g N_VSS_Mn9@4293_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4292 N_OUT9_Mn9@4292_d N_OUT8_Mn9@4292_g N_VSS_Mn9@4292_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4293 N_OUT9_Mp9@4293_d N_OUT8_Mp9@4293_g N_VDD_Mp9@4293_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4292 N_OUT9_Mp9@4292_d N_OUT8_Mp9@4292_g N_VDD_Mp9@4292_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4291 N_OUT9_Mn9@4291_d N_OUT8_Mn9@4291_g N_VSS_Mn9@4291_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4290 N_OUT9_Mn9@4290_d N_OUT8_Mn9@4290_g N_VSS_Mn9@4290_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4291 N_OUT9_Mp9@4291_d N_OUT8_Mp9@4291_g N_VDD_Mp9@4291_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4290 N_OUT9_Mp9@4290_d N_OUT8_Mp9@4290_g N_VDD_Mp9@4290_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4289 N_OUT9_Mn9@4289_d N_OUT8_Mn9@4289_g N_VSS_Mn9@4289_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4288 N_OUT9_Mn9@4288_d N_OUT8_Mn9@4288_g N_VSS_Mn9@4288_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4289 N_OUT9_Mp9@4289_d N_OUT8_Mp9@4289_g N_VDD_Mp9@4289_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4288 N_OUT9_Mp9@4288_d N_OUT8_Mp9@4288_g N_VDD_Mp9@4288_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4287 N_OUT9_Mn9@4287_d N_OUT8_Mn9@4287_g N_VSS_Mn9@4287_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4286 N_OUT9_Mn9@4286_d N_OUT8_Mn9@4286_g N_VSS_Mn9@4286_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4287 N_OUT9_Mp9@4287_d N_OUT8_Mp9@4287_g N_VDD_Mp9@4287_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4286 N_OUT9_Mp9@4286_d N_OUT8_Mp9@4286_g N_VDD_Mp9@4286_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4285 N_OUT9_Mn9@4285_d N_OUT8_Mn9@4285_g N_VSS_Mn9@4285_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4284 N_OUT9_Mn9@4284_d N_OUT8_Mn9@4284_g N_VSS_Mn9@4284_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4285 N_OUT9_Mp9@4285_d N_OUT8_Mp9@4285_g N_VDD_Mp9@4285_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4284 N_OUT9_Mp9@4284_d N_OUT8_Mp9@4284_g N_VDD_Mp9@4284_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4283 N_OUT9_Mn9@4283_d N_OUT8_Mn9@4283_g N_VSS_Mn9@4283_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4282 N_OUT9_Mn9@4282_d N_OUT8_Mn9@4282_g N_VSS_Mn9@4282_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4283 N_OUT9_Mp9@4283_d N_OUT8_Mp9@4283_g N_VDD_Mp9@4283_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4282 N_OUT9_Mp9@4282_d N_OUT8_Mp9@4282_g N_VDD_Mp9@4282_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4281 N_OUT9_Mn9@4281_d N_OUT8_Mn9@4281_g N_VSS_Mn9@4281_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4280 N_OUT9_Mn9@4280_d N_OUT8_Mn9@4280_g N_VSS_Mn9@4280_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4281 N_OUT9_Mp9@4281_d N_OUT8_Mp9@4281_g N_VDD_Mp9@4281_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4280 N_OUT9_Mp9@4280_d N_OUT8_Mp9@4280_g N_VDD_Mp9@4280_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4279 N_OUT9_Mn9@4279_d N_OUT8_Mn9@4279_g N_VSS_Mn9@4279_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4278 N_OUT9_Mn9@4278_d N_OUT8_Mn9@4278_g N_VSS_Mn9@4278_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4279 N_OUT9_Mp9@4279_d N_OUT8_Mp9@4279_g N_VDD_Mp9@4279_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4278 N_OUT9_Mp9@4278_d N_OUT8_Mp9@4278_g N_VDD_Mp9@4278_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4277 N_OUT9_Mn9@4277_d N_OUT8_Mn9@4277_g N_VSS_Mn9@4277_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4276 N_OUT9_Mn9@4276_d N_OUT8_Mn9@4276_g N_VSS_Mn9@4276_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4277 N_OUT9_Mp9@4277_d N_OUT8_Mp9@4277_g N_VDD_Mp9@4277_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4276 N_OUT9_Mp9@4276_d N_OUT8_Mp9@4276_g N_VDD_Mp9@4276_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4275 N_OUT9_Mn9@4275_d N_OUT8_Mn9@4275_g N_VSS_Mn9@4275_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4274 N_OUT9_Mn9@4274_d N_OUT8_Mn9@4274_g N_VSS_Mn9@4274_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4275 N_OUT9_Mp9@4275_d N_OUT8_Mp9@4275_g N_VDD_Mp9@4275_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4274 N_OUT9_Mp9@4274_d N_OUT8_Mp9@4274_g N_VDD_Mp9@4274_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4273 N_OUT9_Mn9@4273_d N_OUT8_Mn9@4273_g N_VSS_Mn9@4273_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4272 N_OUT9_Mn9@4272_d N_OUT8_Mn9@4272_g N_VSS_Mn9@4272_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4273 N_OUT9_Mp9@4273_d N_OUT8_Mp9@4273_g N_VDD_Mp9@4273_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4272 N_OUT9_Mp9@4272_d N_OUT8_Mp9@4272_g N_VDD_Mp9@4272_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4271 N_OUT9_Mn9@4271_d N_OUT8_Mn9@4271_g N_VSS_Mn9@4271_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4270 N_OUT9_Mn9@4270_d N_OUT8_Mn9@4270_g N_VSS_Mn9@4270_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4271 N_OUT9_Mp9@4271_d N_OUT8_Mp9@4271_g N_VDD_Mp9@4271_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4270 N_OUT9_Mp9@4270_d N_OUT8_Mp9@4270_g N_VDD_Mp9@4270_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4269 N_OUT9_Mn9@4269_d N_OUT8_Mn9@4269_g N_VSS_Mn9@4269_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4268 N_OUT9_Mn9@4268_d N_OUT8_Mn9@4268_g N_VSS_Mn9@4268_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4269 N_OUT9_Mp9@4269_d N_OUT8_Mp9@4269_g N_VDD_Mp9@4269_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4268 N_OUT9_Mp9@4268_d N_OUT8_Mp9@4268_g N_VDD_Mp9@4268_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4267 N_OUT9_Mn9@4267_d N_OUT8_Mn9@4267_g N_VSS_Mn9@4267_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4266 N_OUT9_Mn9@4266_d N_OUT8_Mn9@4266_g N_VSS_Mn9@4266_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4267 N_OUT9_Mp9@4267_d N_OUT8_Mp9@4267_g N_VDD_Mp9@4267_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4266 N_OUT9_Mp9@4266_d N_OUT8_Mp9@4266_g N_VDD_Mp9@4266_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4265 N_OUT9_Mn9@4265_d N_OUT8_Mn9@4265_g N_VSS_Mn9@4265_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4264 N_OUT9_Mn9@4264_d N_OUT8_Mn9@4264_g N_VSS_Mn9@4264_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4265 N_OUT9_Mp9@4265_d N_OUT8_Mp9@4265_g N_VDD_Mp9@4265_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4264 N_OUT9_Mp9@4264_d N_OUT8_Mp9@4264_g N_VDD_Mp9@4264_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4263 N_OUT9_Mn9@4263_d N_OUT8_Mn9@4263_g N_VSS_Mn9@4263_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4262 N_OUT9_Mn9@4262_d N_OUT8_Mn9@4262_g N_VSS_Mn9@4262_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4263 N_OUT9_Mp9@4263_d N_OUT8_Mp9@4263_g N_VDD_Mp9@4263_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4262 N_OUT9_Mp9@4262_d N_OUT8_Mp9@4262_g N_VDD_Mp9@4262_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4261 N_OUT9_Mn9@4261_d N_OUT8_Mn9@4261_g N_VSS_Mn9@4261_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4260 N_OUT9_Mn9@4260_d N_OUT8_Mn9@4260_g N_VSS_Mn9@4260_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4261 N_OUT9_Mp9@4261_d N_OUT8_Mp9@4261_g N_VDD_Mp9@4261_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4260 N_OUT9_Mp9@4260_d N_OUT8_Mp9@4260_g N_VDD_Mp9@4260_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4259 N_OUT9_Mn9@4259_d N_OUT8_Mn9@4259_g N_VSS_Mn9@4259_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4258 N_OUT9_Mn9@4258_d N_OUT8_Mn9@4258_g N_VSS_Mn9@4258_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4259 N_OUT9_Mp9@4259_d N_OUT8_Mp9@4259_g N_VDD_Mp9@4259_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4258 N_OUT9_Mp9@4258_d N_OUT8_Mp9@4258_g N_VDD_Mp9@4258_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4257 N_OUT9_Mn9@4257_d N_OUT8_Mn9@4257_g N_VSS_Mn9@4257_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4256 N_OUT9_Mn9@4256_d N_OUT8_Mn9@4256_g N_VSS_Mn9@4256_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4257 N_OUT9_Mp9@4257_d N_OUT8_Mp9@4257_g N_VDD_Mp9@4257_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4256 N_OUT9_Mp9@4256_d N_OUT8_Mp9@4256_g N_VDD_Mp9@4256_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4255 N_OUT9_Mn9@4255_d N_OUT8_Mn9@4255_g N_VSS_Mn9@4255_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4254 N_OUT9_Mn9@4254_d N_OUT8_Mn9@4254_g N_VSS_Mn9@4254_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4255 N_OUT9_Mp9@4255_d N_OUT8_Mp9@4255_g N_VDD_Mp9@4255_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4254 N_OUT9_Mp9@4254_d N_OUT8_Mp9@4254_g N_VDD_Mp9@4254_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4253 N_OUT9_Mn9@4253_d N_OUT8_Mn9@4253_g N_VSS_Mn9@4253_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4252 N_OUT9_Mn9@4252_d N_OUT8_Mn9@4252_g N_VSS_Mn9@4252_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4253 N_OUT9_Mp9@4253_d N_OUT8_Mp9@4253_g N_VDD_Mp9@4253_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4252 N_OUT9_Mp9@4252_d N_OUT8_Mp9@4252_g N_VDD_Mp9@4252_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4251 N_OUT9_Mn9@4251_d N_OUT8_Mn9@4251_g N_VSS_Mn9@4251_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4250 N_OUT9_Mn9@4250_d N_OUT8_Mn9@4250_g N_VSS_Mn9@4250_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4251 N_OUT9_Mp9@4251_d N_OUT8_Mp9@4251_g N_VDD_Mp9@4251_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4250 N_OUT9_Mp9@4250_d N_OUT8_Mp9@4250_g N_VDD_Mp9@4250_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4249 N_OUT9_Mn9@4249_d N_OUT8_Mn9@4249_g N_VSS_Mn9@4249_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4248 N_OUT9_Mn9@4248_d N_OUT8_Mn9@4248_g N_VSS_Mn9@4248_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4249 N_OUT9_Mp9@4249_d N_OUT8_Mp9@4249_g N_VDD_Mp9@4249_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4248 N_OUT9_Mp9@4248_d N_OUT8_Mp9@4248_g N_VDD_Mp9@4248_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4247 N_OUT9_Mn9@4247_d N_OUT8_Mn9@4247_g N_VSS_Mn9@4247_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4246 N_OUT9_Mn9@4246_d N_OUT8_Mn9@4246_g N_VSS_Mn9@4246_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4247 N_OUT9_Mp9@4247_d N_OUT8_Mp9@4247_g N_VDD_Mp9@4247_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4246 N_OUT9_Mp9@4246_d N_OUT8_Mp9@4246_g N_VDD_Mp9@4246_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4245 N_OUT9_Mn9@4245_d N_OUT8_Mn9@4245_g N_VSS_Mn9@4245_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4244 N_OUT9_Mn9@4244_d N_OUT8_Mn9@4244_g N_VSS_Mn9@4244_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4245 N_OUT9_Mp9@4245_d N_OUT8_Mp9@4245_g N_VDD_Mp9@4245_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4244 N_OUT9_Mp9@4244_d N_OUT8_Mp9@4244_g N_VDD_Mp9@4244_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4243 N_OUT9_Mn9@4243_d N_OUT8_Mn9@4243_g N_VSS_Mn9@4243_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4242 N_OUT9_Mn9@4242_d N_OUT8_Mn9@4242_g N_VSS_Mn9@4242_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4243 N_OUT9_Mp9@4243_d N_OUT8_Mp9@4243_g N_VDD_Mp9@4243_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4242 N_OUT9_Mp9@4242_d N_OUT8_Mp9@4242_g N_VDD_Mp9@4242_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4241 N_OUT9_Mn9@4241_d N_OUT8_Mn9@4241_g N_VSS_Mn9@4241_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4240 N_OUT9_Mn9@4240_d N_OUT8_Mn9@4240_g N_VSS_Mn9@4240_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4241 N_OUT9_Mp9@4241_d N_OUT8_Mp9@4241_g N_VDD_Mp9@4241_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4240 N_OUT9_Mp9@4240_d N_OUT8_Mp9@4240_g N_VDD_Mp9@4240_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4239 N_OUT9_Mn9@4239_d N_OUT8_Mn9@4239_g N_VSS_Mn9@4239_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4238 N_OUT9_Mn9@4238_d N_OUT8_Mn9@4238_g N_VSS_Mn9@4238_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4239 N_OUT9_Mp9@4239_d N_OUT8_Mp9@4239_g N_VDD_Mp9@4239_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4238 N_OUT9_Mp9@4238_d N_OUT8_Mp9@4238_g N_VDD_Mp9@4238_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4237 N_OUT9_Mn9@4237_d N_OUT8_Mn9@4237_g N_VSS_Mn9@4237_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4236 N_OUT9_Mn9@4236_d N_OUT8_Mn9@4236_g N_VSS_Mn9@4236_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4237 N_OUT9_Mp9@4237_d N_OUT8_Mp9@4237_g N_VDD_Mp9@4237_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4236 N_OUT9_Mp9@4236_d N_OUT8_Mp9@4236_g N_VDD_Mp9@4236_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4235 N_OUT9_Mn9@4235_d N_OUT8_Mn9@4235_g N_VSS_Mn9@4235_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4234 N_OUT9_Mn9@4234_d N_OUT8_Mn9@4234_g N_VSS_Mn9@4234_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4235 N_OUT9_Mp9@4235_d N_OUT8_Mp9@4235_g N_VDD_Mp9@4235_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4234 N_OUT9_Mp9@4234_d N_OUT8_Mp9@4234_g N_VDD_Mp9@4234_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4233 N_OUT9_Mn9@4233_d N_OUT8_Mn9@4233_g N_VSS_Mn9@4233_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4232 N_OUT9_Mn9@4232_d N_OUT8_Mn9@4232_g N_VSS_Mn9@4232_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4233 N_OUT9_Mp9@4233_d N_OUT8_Mp9@4233_g N_VDD_Mp9@4233_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4232 N_OUT9_Mp9@4232_d N_OUT8_Mp9@4232_g N_VDD_Mp9@4232_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4231 N_OUT9_Mn9@4231_d N_OUT8_Mn9@4231_g N_VSS_Mn9@4231_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4230 N_OUT9_Mn9@4230_d N_OUT8_Mn9@4230_g N_VSS_Mn9@4230_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4231 N_OUT9_Mp9@4231_d N_OUT8_Mp9@4231_g N_VDD_Mp9@4231_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4230 N_OUT9_Mp9@4230_d N_OUT8_Mp9@4230_g N_VDD_Mp9@4230_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4229 N_OUT9_Mn9@4229_d N_OUT8_Mn9@4229_g N_VSS_Mn9@4229_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4228 N_OUT9_Mn9@4228_d N_OUT8_Mn9@4228_g N_VSS_Mn9@4228_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4229 N_OUT9_Mp9@4229_d N_OUT8_Mp9@4229_g N_VDD_Mp9@4229_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4228 N_OUT9_Mp9@4228_d N_OUT8_Mp9@4228_g N_VDD_Mp9@4228_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4227 N_OUT9_Mn9@4227_d N_OUT8_Mn9@4227_g N_VSS_Mn9@4227_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4226 N_OUT9_Mn9@4226_d N_OUT8_Mn9@4226_g N_VSS_Mn9@4226_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4227 N_OUT9_Mp9@4227_d N_OUT8_Mp9@4227_g N_VDD_Mp9@4227_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4226 N_OUT9_Mp9@4226_d N_OUT8_Mp9@4226_g N_VDD_Mp9@4226_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4225 N_OUT9_Mn9@4225_d N_OUT8_Mn9@4225_g N_VSS_Mn9@4225_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4224 N_OUT9_Mn9@4224_d N_OUT8_Mn9@4224_g N_VSS_Mn9@4224_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4225 N_OUT9_Mp9@4225_d N_OUT8_Mp9@4225_g N_VDD_Mp9@4225_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4224 N_OUT9_Mp9@4224_d N_OUT8_Mp9@4224_g N_VDD_Mp9@4224_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4223 N_OUT9_Mn9@4223_d N_OUT8_Mn9@4223_g N_VSS_Mn9@4223_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4222 N_OUT9_Mn9@4222_d N_OUT8_Mn9@4222_g N_VSS_Mn9@4222_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4223 N_OUT9_Mp9@4223_d N_OUT8_Mp9@4223_g N_VDD_Mp9@4223_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4222 N_OUT9_Mp9@4222_d N_OUT8_Mp9@4222_g N_VDD_Mp9@4222_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4221 N_OUT9_Mn9@4221_d N_OUT8_Mn9@4221_g N_VSS_Mn9@4221_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4220 N_OUT9_Mn9@4220_d N_OUT8_Mn9@4220_g N_VSS_Mn9@4220_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4221 N_OUT9_Mp9@4221_d N_OUT8_Mp9@4221_g N_VDD_Mp9@4221_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4220 N_OUT9_Mp9@4220_d N_OUT8_Mp9@4220_g N_VDD_Mp9@4220_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4219 N_OUT9_Mn9@4219_d N_OUT8_Mn9@4219_g N_VSS_Mn9@4219_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4218 N_OUT9_Mn9@4218_d N_OUT8_Mn9@4218_g N_VSS_Mn9@4218_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4219 N_OUT9_Mp9@4219_d N_OUT8_Mp9@4219_g N_VDD_Mp9@4219_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4218 N_OUT9_Mp9@4218_d N_OUT8_Mp9@4218_g N_VDD_Mp9@4218_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4217 N_OUT9_Mn9@4217_d N_OUT8_Mn9@4217_g N_VSS_Mn9@4217_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4216 N_OUT9_Mn9@4216_d N_OUT8_Mn9@4216_g N_VSS_Mn9@4216_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4217 N_OUT9_Mp9@4217_d N_OUT8_Mp9@4217_g N_VDD_Mp9@4217_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4216 N_OUT9_Mp9@4216_d N_OUT8_Mp9@4216_g N_VDD_Mp9@4216_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4215 N_OUT9_Mn9@4215_d N_OUT8_Mn9@4215_g N_VSS_Mn9@4215_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4214 N_OUT9_Mn9@4214_d N_OUT8_Mn9@4214_g N_VSS_Mn9@4214_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4215 N_OUT9_Mp9@4215_d N_OUT8_Mp9@4215_g N_VDD_Mp9@4215_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4214 N_OUT9_Mp9@4214_d N_OUT8_Mp9@4214_g N_VDD_Mp9@4214_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4213 N_OUT9_Mn9@4213_d N_OUT8_Mn9@4213_g N_VSS_Mn9@4213_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4212 N_OUT9_Mn9@4212_d N_OUT8_Mn9@4212_g N_VSS_Mn9@4212_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4213 N_OUT9_Mp9@4213_d N_OUT8_Mp9@4213_g N_VDD_Mp9@4213_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4212 N_OUT9_Mp9@4212_d N_OUT8_Mp9@4212_g N_VDD_Mp9@4212_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4211 N_OUT9_Mn9@4211_d N_OUT8_Mn9@4211_g N_VSS_Mn9@4211_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4210 N_OUT9_Mn9@4210_d N_OUT8_Mn9@4210_g N_VSS_Mn9@4210_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4211 N_OUT9_Mp9@4211_d N_OUT8_Mp9@4211_g N_VDD_Mp9@4211_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4210 N_OUT9_Mp9@4210_d N_OUT8_Mp9@4210_g N_VDD_Mp9@4210_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4209 N_OUT9_Mn9@4209_d N_OUT8_Mn9@4209_g N_VSS_Mn9@4209_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4208 N_OUT9_Mn9@4208_d N_OUT8_Mn9@4208_g N_VSS_Mn9@4208_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4209 N_OUT9_Mp9@4209_d N_OUT8_Mp9@4209_g N_VDD_Mp9@4209_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4208 N_OUT9_Mp9@4208_d N_OUT8_Mp9@4208_g N_VDD_Mp9@4208_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4207 N_OUT9_Mn9@4207_d N_OUT8_Mn9@4207_g N_VSS_Mn9@4207_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4206 N_OUT9_Mn9@4206_d N_OUT8_Mn9@4206_g N_VSS_Mn9@4206_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4207 N_OUT9_Mp9@4207_d N_OUT8_Mp9@4207_g N_VDD_Mp9@4207_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4206 N_OUT9_Mp9@4206_d N_OUT8_Mp9@4206_g N_VDD_Mp9@4206_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4205 N_OUT9_Mn9@4205_d N_OUT8_Mn9@4205_g N_VSS_Mn9@4205_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4204 N_OUT9_Mn9@4204_d N_OUT8_Mn9@4204_g N_VSS_Mn9@4204_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4205 N_OUT9_Mp9@4205_d N_OUT8_Mp9@4205_g N_VDD_Mp9@4205_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4204 N_OUT9_Mp9@4204_d N_OUT8_Mp9@4204_g N_VDD_Mp9@4204_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4203 N_OUT9_Mn9@4203_d N_OUT8_Mn9@4203_g N_VSS_Mn9@4203_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4202 N_OUT9_Mn9@4202_d N_OUT8_Mn9@4202_g N_VSS_Mn9@4202_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4203 N_OUT9_Mp9@4203_d N_OUT8_Mp9@4203_g N_VDD_Mp9@4203_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4202 N_OUT9_Mp9@4202_d N_OUT8_Mp9@4202_g N_VDD_Mp9@4202_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4201 N_OUT9_Mn9@4201_d N_OUT8_Mn9@4201_g N_VSS_Mn9@4201_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4200 N_OUT9_Mn9@4200_d N_OUT8_Mn9@4200_g N_VSS_Mn9@4200_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4201 N_OUT9_Mp9@4201_d N_OUT8_Mp9@4201_g N_VDD_Mp9@4201_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4200 N_OUT9_Mp9@4200_d N_OUT8_Mp9@4200_g N_VDD_Mp9@4200_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4199 N_OUT9_Mn9@4199_d N_OUT8_Mn9@4199_g N_VSS_Mn9@4199_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4198 N_OUT9_Mn9@4198_d N_OUT8_Mn9@4198_g N_VSS_Mn9@4198_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4199 N_OUT9_Mp9@4199_d N_OUT8_Mp9@4199_g N_VDD_Mp9@4199_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4198 N_OUT9_Mp9@4198_d N_OUT8_Mp9@4198_g N_VDD_Mp9@4198_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4197 N_OUT9_Mn9@4197_d N_OUT8_Mn9@4197_g N_VSS_Mn9@4197_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4196 N_OUT9_Mn9@4196_d N_OUT8_Mn9@4196_g N_VSS_Mn9@4196_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4197 N_OUT9_Mp9@4197_d N_OUT8_Mp9@4197_g N_VDD_Mp9@4197_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4196 N_OUT9_Mp9@4196_d N_OUT8_Mp9@4196_g N_VDD_Mp9@4196_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4195 N_OUT9_Mn9@4195_d N_OUT8_Mn9@4195_g N_VSS_Mn9@4195_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4194 N_OUT9_Mn9@4194_d N_OUT8_Mn9@4194_g N_VSS_Mn9@4194_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4195 N_OUT9_Mp9@4195_d N_OUT8_Mp9@4195_g N_VDD_Mp9@4195_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4194 N_OUT9_Mp9@4194_d N_OUT8_Mp9@4194_g N_VDD_Mp9@4194_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4193 N_OUT9_Mn9@4193_d N_OUT8_Mn9@4193_g N_VSS_Mn9@4193_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4192 N_OUT9_Mn9@4192_d N_OUT8_Mn9@4192_g N_VSS_Mn9@4192_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4193 N_OUT9_Mp9@4193_d N_OUT8_Mp9@4193_g N_VDD_Mp9@4193_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4192 N_OUT9_Mp9@4192_d N_OUT8_Mp9@4192_g N_VDD_Mp9@4192_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4191 N_OUT9_Mn9@4191_d N_OUT8_Mn9@4191_g N_VSS_Mn9@4191_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4190 N_OUT9_Mn9@4190_d N_OUT8_Mn9@4190_g N_VSS_Mn9@4190_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4191 N_OUT9_Mp9@4191_d N_OUT8_Mp9@4191_g N_VDD_Mp9@4191_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4190 N_OUT9_Mp9@4190_d N_OUT8_Mp9@4190_g N_VDD_Mp9@4190_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4189 N_OUT9_Mn9@4189_d N_OUT8_Mn9@4189_g N_VSS_Mn9@4189_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4188 N_OUT9_Mn9@4188_d N_OUT8_Mn9@4188_g N_VSS_Mn9@4188_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4189 N_OUT9_Mp9@4189_d N_OUT8_Mp9@4189_g N_VDD_Mp9@4189_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4188 N_OUT9_Mp9@4188_d N_OUT8_Mp9@4188_g N_VDD_Mp9@4188_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4187 N_OUT9_Mn9@4187_d N_OUT8_Mn9@4187_g N_VSS_Mn9@4187_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4186 N_OUT9_Mn9@4186_d N_OUT8_Mn9@4186_g N_VSS_Mn9@4186_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4187 N_OUT9_Mp9@4187_d N_OUT8_Mp9@4187_g N_VDD_Mp9@4187_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4186 N_OUT9_Mp9@4186_d N_OUT8_Mp9@4186_g N_VDD_Mp9@4186_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4185 N_OUT9_Mn9@4185_d N_OUT8_Mn9@4185_g N_VSS_Mn9@4185_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4184 N_OUT9_Mn9@4184_d N_OUT8_Mn9@4184_g N_VSS_Mn9@4184_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4185 N_OUT9_Mp9@4185_d N_OUT8_Mp9@4185_g N_VDD_Mp9@4185_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4184 N_OUT9_Mp9@4184_d N_OUT8_Mp9@4184_g N_VDD_Mp9@4184_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4183 N_OUT9_Mn9@4183_d N_OUT8_Mn9@4183_g N_VSS_Mn9@4183_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4182 N_OUT9_Mn9@4182_d N_OUT8_Mn9@4182_g N_VSS_Mn9@4182_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4183 N_OUT9_Mp9@4183_d N_OUT8_Mp9@4183_g N_VDD_Mp9@4183_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4182 N_OUT9_Mp9@4182_d N_OUT8_Mp9@4182_g N_VDD_Mp9@4182_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4181 N_OUT9_Mn9@4181_d N_OUT8_Mn9@4181_g N_VSS_Mn9@4181_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4180 N_OUT9_Mn9@4180_d N_OUT8_Mn9@4180_g N_VSS_Mn9@4180_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4181 N_OUT9_Mp9@4181_d N_OUT8_Mp9@4181_g N_VDD_Mp9@4181_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4180 N_OUT9_Mp9@4180_d N_OUT8_Mp9@4180_g N_VDD_Mp9@4180_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4179 N_OUT9_Mn9@4179_d N_OUT8_Mn9@4179_g N_VSS_Mn9@4179_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4178 N_OUT9_Mn9@4178_d N_OUT8_Mn9@4178_g N_VSS_Mn9@4178_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4179 N_OUT9_Mp9@4179_d N_OUT8_Mp9@4179_g N_VDD_Mp9@4179_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4178 N_OUT9_Mp9@4178_d N_OUT8_Mp9@4178_g N_VDD_Mp9@4178_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4177 N_OUT9_Mn9@4177_d N_OUT8_Mn9@4177_g N_VSS_Mn9@4177_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4176 N_OUT9_Mn9@4176_d N_OUT8_Mn9@4176_g N_VSS_Mn9@4176_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4177 N_OUT9_Mp9@4177_d N_OUT8_Mp9@4177_g N_VDD_Mp9@4177_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4176 N_OUT9_Mp9@4176_d N_OUT8_Mp9@4176_g N_VDD_Mp9@4176_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4175 N_OUT9_Mn9@4175_d N_OUT8_Mn9@4175_g N_VSS_Mn9@4175_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4174 N_OUT9_Mn9@4174_d N_OUT8_Mn9@4174_g N_VSS_Mn9@4174_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4175 N_OUT9_Mp9@4175_d N_OUT8_Mp9@4175_g N_VDD_Mp9@4175_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4174 N_OUT9_Mp9@4174_d N_OUT8_Mp9@4174_g N_VDD_Mp9@4174_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4173 N_OUT9_Mn9@4173_d N_OUT8_Mn9@4173_g N_VSS_Mn9@4173_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4172 N_OUT9_Mn9@4172_d N_OUT8_Mn9@4172_g N_VSS_Mn9@4172_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4173 N_OUT9_Mp9@4173_d N_OUT8_Mp9@4173_g N_VDD_Mp9@4173_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4172 N_OUT9_Mp9@4172_d N_OUT8_Mp9@4172_g N_VDD_Mp9@4172_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4171 N_OUT9_Mn9@4171_d N_OUT8_Mn9@4171_g N_VSS_Mn9@4171_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4170 N_OUT9_Mn9@4170_d N_OUT8_Mn9@4170_g N_VSS_Mn9@4170_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4171 N_OUT9_Mp9@4171_d N_OUT8_Mp9@4171_g N_VDD_Mp9@4171_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4170 N_OUT9_Mp9@4170_d N_OUT8_Mp9@4170_g N_VDD_Mp9@4170_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4169 N_OUT9_Mn9@4169_d N_OUT8_Mn9@4169_g N_VSS_Mn9@4169_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4168 N_OUT9_Mn9@4168_d N_OUT8_Mn9@4168_g N_VSS_Mn9@4168_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4169 N_OUT9_Mp9@4169_d N_OUT8_Mp9@4169_g N_VDD_Mp9@4169_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4168 N_OUT9_Mp9@4168_d N_OUT8_Mp9@4168_g N_VDD_Mp9@4168_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4167 N_OUT9_Mn9@4167_d N_OUT8_Mn9@4167_g N_VSS_Mn9@4167_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4166 N_OUT9_Mn9@4166_d N_OUT8_Mn9@4166_g N_VSS_Mn9@4166_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4167 N_OUT9_Mp9@4167_d N_OUT8_Mp9@4167_g N_VDD_Mp9@4167_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4166 N_OUT9_Mp9@4166_d N_OUT8_Mp9@4166_g N_VDD_Mp9@4166_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4165 N_OUT9_Mn9@4165_d N_OUT8_Mn9@4165_g N_VSS_Mn9@4165_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4164 N_OUT9_Mn9@4164_d N_OUT8_Mn9@4164_g N_VSS_Mn9@4164_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4165 N_OUT9_Mp9@4165_d N_OUT8_Mp9@4165_g N_VDD_Mp9@4165_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4164 N_OUT9_Mp9@4164_d N_OUT8_Mp9@4164_g N_VDD_Mp9@4164_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4163 N_OUT9_Mn9@4163_d N_OUT8_Mn9@4163_g N_VSS_Mn9@4163_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4162 N_OUT9_Mn9@4162_d N_OUT8_Mn9@4162_g N_VSS_Mn9@4162_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4163 N_OUT9_Mp9@4163_d N_OUT8_Mp9@4163_g N_VDD_Mp9@4163_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4162 N_OUT9_Mp9@4162_d N_OUT8_Mp9@4162_g N_VDD_Mp9@4162_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4161 N_OUT9_Mn9@4161_d N_OUT8_Mn9@4161_g N_VSS_Mn9@4161_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4160 N_OUT9_Mn9@4160_d N_OUT8_Mn9@4160_g N_VSS_Mn9@4160_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4161 N_OUT9_Mp9@4161_d N_OUT8_Mp9@4161_g N_VDD_Mp9@4161_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4160 N_OUT9_Mp9@4160_d N_OUT8_Mp9@4160_g N_VDD_Mp9@4160_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4159 N_OUT9_Mn9@4159_d N_OUT8_Mn9@4159_g N_VSS_Mn9@4159_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4158 N_OUT9_Mn9@4158_d N_OUT8_Mn9@4158_g N_VSS_Mn9@4158_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4159 N_OUT9_Mp9@4159_d N_OUT8_Mp9@4159_g N_VDD_Mp9@4159_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4158 N_OUT9_Mp9@4158_d N_OUT8_Mp9@4158_g N_VDD_Mp9@4158_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4157 N_OUT9_Mn9@4157_d N_OUT8_Mn9@4157_g N_VSS_Mn9@4157_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4156 N_OUT9_Mn9@4156_d N_OUT8_Mn9@4156_g N_VSS_Mn9@4156_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4157 N_OUT9_Mp9@4157_d N_OUT8_Mp9@4157_g N_VDD_Mp9@4157_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4156 N_OUT9_Mp9@4156_d N_OUT8_Mp9@4156_g N_VDD_Mp9@4156_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4155 N_OUT9_Mn9@4155_d N_OUT8_Mn9@4155_g N_VSS_Mn9@4155_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4154 N_OUT9_Mn9@4154_d N_OUT8_Mn9@4154_g N_VSS_Mn9@4154_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4155 N_OUT9_Mp9@4155_d N_OUT8_Mp9@4155_g N_VDD_Mp9@4155_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4154 N_OUT9_Mp9@4154_d N_OUT8_Mp9@4154_g N_VDD_Mp9@4154_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4153 N_OUT9_Mn9@4153_d N_OUT8_Mn9@4153_g N_VSS_Mn9@4153_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4152 N_OUT9_Mn9@4152_d N_OUT8_Mn9@4152_g N_VSS_Mn9@4152_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4153 N_OUT9_Mp9@4153_d N_OUT8_Mp9@4153_g N_VDD_Mp9@4153_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4152 N_OUT9_Mp9@4152_d N_OUT8_Mp9@4152_g N_VDD_Mp9@4152_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4151 N_OUT9_Mn9@4151_d N_OUT8_Mn9@4151_g N_VSS_Mn9@4151_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4150 N_OUT9_Mn9@4150_d N_OUT8_Mn9@4150_g N_VSS_Mn9@4150_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4151 N_OUT9_Mp9@4151_d N_OUT8_Mp9@4151_g N_VDD_Mp9@4151_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4150 N_OUT9_Mp9@4150_d N_OUT8_Mp9@4150_g N_VDD_Mp9@4150_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4149 N_OUT9_Mn9@4149_d N_OUT8_Mn9@4149_g N_VSS_Mn9@4149_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4148 N_OUT9_Mn9@4148_d N_OUT8_Mn9@4148_g N_VSS_Mn9@4148_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4149 N_OUT9_Mp9@4149_d N_OUT8_Mp9@4149_g N_VDD_Mp9@4149_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4148 N_OUT9_Mp9@4148_d N_OUT8_Mp9@4148_g N_VDD_Mp9@4148_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4147 N_OUT9_Mn9@4147_d N_OUT8_Mn9@4147_g N_VSS_Mn9@4147_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4146 N_OUT9_Mn9@4146_d N_OUT8_Mn9@4146_g N_VSS_Mn9@4146_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4147 N_OUT9_Mp9@4147_d N_OUT8_Mp9@4147_g N_VDD_Mp9@4147_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4146 N_OUT9_Mp9@4146_d N_OUT8_Mp9@4146_g N_VDD_Mp9@4146_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4145 N_OUT9_Mn9@4145_d N_OUT8_Mn9@4145_g N_VSS_Mn9@4145_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4144 N_OUT9_Mn9@4144_d N_OUT8_Mn9@4144_g N_VSS_Mn9@4144_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4145 N_OUT9_Mp9@4145_d N_OUT8_Mp9@4145_g N_VDD_Mp9@4145_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4144 N_OUT9_Mp9@4144_d N_OUT8_Mp9@4144_g N_VDD_Mp9@4144_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4143 N_OUT9_Mn9@4143_d N_OUT8_Mn9@4143_g N_VSS_Mn9@4143_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4142 N_OUT9_Mn9@4142_d N_OUT8_Mn9@4142_g N_VSS_Mn9@4142_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4143 N_OUT9_Mp9@4143_d N_OUT8_Mp9@4143_g N_VDD_Mp9@4143_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4142 N_OUT9_Mp9@4142_d N_OUT8_Mp9@4142_g N_VDD_Mp9@4142_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4141 N_OUT9_Mn9@4141_d N_OUT8_Mn9@4141_g N_VSS_Mn9@4141_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4140 N_OUT9_Mn9@4140_d N_OUT8_Mn9@4140_g N_VSS_Mn9@4140_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4141 N_OUT9_Mp9@4141_d N_OUT8_Mp9@4141_g N_VDD_Mp9@4141_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4140 N_OUT9_Mp9@4140_d N_OUT8_Mp9@4140_g N_VDD_Mp9@4140_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4139 N_OUT9_Mn9@4139_d N_OUT8_Mn9@4139_g N_VSS_Mn9@4139_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4138 N_OUT9_Mn9@4138_d N_OUT8_Mn9@4138_g N_VSS_Mn9@4138_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4139 N_OUT9_Mp9@4139_d N_OUT8_Mp9@4139_g N_VDD_Mp9@4139_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4138 N_OUT9_Mp9@4138_d N_OUT8_Mp9@4138_g N_VDD_Mp9@4138_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4137 N_OUT9_Mn9@4137_d N_OUT8_Mn9@4137_g N_VSS_Mn9@4137_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4136 N_OUT9_Mn9@4136_d N_OUT8_Mn9@4136_g N_VSS_Mn9@4136_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4137 N_OUT9_Mp9@4137_d N_OUT8_Mp9@4137_g N_VDD_Mp9@4137_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4136 N_OUT9_Mp9@4136_d N_OUT8_Mp9@4136_g N_VDD_Mp9@4136_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4135 N_OUT9_Mn9@4135_d N_OUT8_Mn9@4135_g N_VSS_Mn9@4135_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4134 N_OUT9_Mn9@4134_d N_OUT8_Mn9@4134_g N_VSS_Mn9@4134_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4135 N_OUT9_Mp9@4135_d N_OUT8_Mp9@4135_g N_VDD_Mp9@4135_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4134 N_OUT9_Mp9@4134_d N_OUT8_Mp9@4134_g N_VDD_Mp9@4134_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4133 N_OUT9_Mn9@4133_d N_OUT8_Mn9@4133_g N_VSS_Mn9@4133_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4132 N_OUT9_Mn9@4132_d N_OUT8_Mn9@4132_g N_VSS_Mn9@4132_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4133 N_OUT9_Mp9@4133_d N_OUT8_Mp9@4133_g N_VDD_Mp9@4133_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4132 N_OUT9_Mp9@4132_d N_OUT8_Mp9@4132_g N_VDD_Mp9@4132_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4131 N_OUT9_Mn9@4131_d N_OUT8_Mn9@4131_g N_VSS_Mn9@4131_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4130 N_OUT9_Mn9@4130_d N_OUT8_Mn9@4130_g N_VSS_Mn9@4130_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4131 N_OUT9_Mp9@4131_d N_OUT8_Mp9@4131_g N_VDD_Mp9@4131_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4130 N_OUT9_Mp9@4130_d N_OUT8_Mp9@4130_g N_VDD_Mp9@4130_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4129 N_OUT9_Mn9@4129_d N_OUT8_Mn9@4129_g N_VSS_Mn9@4129_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4128 N_OUT9_Mn9@4128_d N_OUT8_Mn9@4128_g N_VSS_Mn9@4128_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4129 N_OUT9_Mp9@4129_d N_OUT8_Mp9@4129_g N_VDD_Mp9@4129_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4128 N_OUT9_Mp9@4128_d N_OUT8_Mp9@4128_g N_VDD_Mp9@4128_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4127 N_OUT9_Mn9@4127_d N_OUT8_Mn9@4127_g N_VSS_Mn9@4127_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4126 N_OUT9_Mn9@4126_d N_OUT8_Mn9@4126_g N_VSS_Mn9@4126_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4127 N_OUT9_Mp9@4127_d N_OUT8_Mp9@4127_g N_VDD_Mp9@4127_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4126 N_OUT9_Mp9@4126_d N_OUT8_Mp9@4126_g N_VDD_Mp9@4126_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4125 N_OUT9_Mn9@4125_d N_OUT8_Mn9@4125_g N_VSS_Mn9@4125_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4124 N_OUT9_Mn9@4124_d N_OUT8_Mn9@4124_g N_VSS_Mn9@4124_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4125 N_OUT9_Mp9@4125_d N_OUT8_Mp9@4125_g N_VDD_Mp9@4125_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4124 N_OUT9_Mp9@4124_d N_OUT8_Mp9@4124_g N_VDD_Mp9@4124_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4123 N_OUT9_Mn9@4123_d N_OUT8_Mn9@4123_g N_VSS_Mn9@4123_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4122 N_OUT9_Mn9@4122_d N_OUT8_Mn9@4122_g N_VSS_Mn9@4122_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4123 N_OUT9_Mp9@4123_d N_OUT8_Mp9@4123_g N_VDD_Mp9@4123_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4122 N_OUT9_Mp9@4122_d N_OUT8_Mp9@4122_g N_VDD_Mp9@4122_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4121 N_OUT9_Mn9@4121_d N_OUT8_Mn9@4121_g N_VSS_Mn9@4121_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4120 N_OUT9_Mn9@4120_d N_OUT8_Mn9@4120_g N_VSS_Mn9@4120_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4121 N_OUT9_Mp9@4121_d N_OUT8_Mp9@4121_g N_VDD_Mp9@4121_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4120 N_OUT9_Mp9@4120_d N_OUT8_Mp9@4120_g N_VDD_Mp9@4120_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4119 N_OUT9_Mn9@4119_d N_OUT8_Mn9@4119_g N_VSS_Mn9@4119_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4118 N_OUT9_Mn9@4118_d N_OUT8_Mn9@4118_g N_VSS_Mn9@4118_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4119 N_OUT9_Mp9@4119_d N_OUT8_Mp9@4119_g N_VDD_Mp9@4119_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4118 N_OUT9_Mp9@4118_d N_OUT8_Mp9@4118_g N_VDD_Mp9@4118_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4117 N_OUT9_Mn9@4117_d N_OUT8_Mn9@4117_g N_VSS_Mn9@4117_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4116 N_OUT9_Mn9@4116_d N_OUT8_Mn9@4116_g N_VSS_Mn9@4116_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4117 N_OUT9_Mp9@4117_d N_OUT8_Mp9@4117_g N_VDD_Mp9@4117_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4116 N_OUT9_Mp9@4116_d N_OUT8_Mp9@4116_g N_VDD_Mp9@4116_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4115 N_OUT9_Mn9@4115_d N_OUT8_Mn9@4115_g N_VSS_Mn9@4115_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4114 N_OUT9_Mn9@4114_d N_OUT8_Mn9@4114_g N_VSS_Mn9@4114_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4115 N_OUT9_Mp9@4115_d N_OUT8_Mp9@4115_g N_VDD_Mp9@4115_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4114 N_OUT9_Mp9@4114_d N_OUT8_Mp9@4114_g N_VDD_Mp9@4114_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4113 N_OUT9_Mn9@4113_d N_OUT8_Mn9@4113_g N_VSS_Mn9@4113_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4112 N_OUT9_Mn9@4112_d N_OUT8_Mn9@4112_g N_VSS_Mn9@4112_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4113 N_OUT9_Mp9@4113_d N_OUT8_Mp9@4113_g N_VDD_Mp9@4113_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4112 N_OUT9_Mp9@4112_d N_OUT8_Mp9@4112_g N_VDD_Mp9@4112_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4111 N_OUT9_Mn9@4111_d N_OUT8_Mn9@4111_g N_VSS_Mn9@4111_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4110 N_OUT9_Mn9@4110_d N_OUT8_Mn9@4110_g N_VSS_Mn9@4110_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4111 N_OUT9_Mp9@4111_d N_OUT8_Mp9@4111_g N_VDD_Mp9@4111_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4110 N_OUT9_Mp9@4110_d N_OUT8_Mp9@4110_g N_VDD_Mp9@4110_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4109 N_OUT9_Mn9@4109_d N_OUT8_Mn9@4109_g N_VSS_Mn9@4109_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4108 N_OUT9_Mn9@4108_d N_OUT8_Mn9@4108_g N_VSS_Mn9@4108_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4109 N_OUT9_Mp9@4109_d N_OUT8_Mp9@4109_g N_VDD_Mp9@4109_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4108 N_OUT9_Mp9@4108_d N_OUT8_Mp9@4108_g N_VDD_Mp9@4108_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4107 N_OUT9_Mn9@4107_d N_OUT8_Mn9@4107_g N_VSS_Mn9@4107_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4106 N_OUT9_Mn9@4106_d N_OUT8_Mn9@4106_g N_VSS_Mn9@4106_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4107 N_OUT9_Mp9@4107_d N_OUT8_Mp9@4107_g N_VDD_Mp9@4107_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4106 N_OUT9_Mp9@4106_d N_OUT8_Mp9@4106_g N_VDD_Mp9@4106_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4105 N_OUT9_Mn9@4105_d N_OUT8_Mn9@4105_g N_VSS_Mn9@4105_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4104 N_OUT9_Mn9@4104_d N_OUT8_Mn9@4104_g N_VSS_Mn9@4104_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4105 N_OUT9_Mp9@4105_d N_OUT8_Mp9@4105_g N_VDD_Mp9@4105_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4104 N_OUT9_Mp9@4104_d N_OUT8_Mp9@4104_g N_VDD_Mp9@4104_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4103 N_OUT9_Mn9@4103_d N_OUT8_Mn9@4103_g N_VSS_Mn9@4103_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4102 N_OUT9_Mn9@4102_d N_OUT8_Mn9@4102_g N_VSS_Mn9@4102_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4103 N_OUT9_Mp9@4103_d N_OUT8_Mp9@4103_g N_VDD_Mp9@4103_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4102 N_OUT9_Mp9@4102_d N_OUT8_Mp9@4102_g N_VDD_Mp9@4102_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4101 N_OUT9_Mn9@4101_d N_OUT8_Mn9@4101_g N_VSS_Mn9@4101_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4100 N_OUT9_Mn9@4100_d N_OUT8_Mn9@4100_g N_VSS_Mn9@4100_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4101 N_OUT9_Mp9@4101_d N_OUT8_Mp9@4101_g N_VDD_Mp9@4101_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4100 N_OUT9_Mp9@4100_d N_OUT8_Mp9@4100_g N_VDD_Mp9@4100_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4099 N_OUT9_Mn9@4099_d N_OUT8_Mn9@4099_g N_VSS_Mn9@4099_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4098 N_OUT9_Mn9@4098_d N_OUT8_Mn9@4098_g N_VSS_Mn9@4098_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4099 N_OUT9_Mp9@4099_d N_OUT8_Mp9@4099_g N_VDD_Mp9@4099_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4098 N_OUT9_Mp9@4098_d N_OUT8_Mp9@4098_g N_VDD_Mp9@4098_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1025 N_OUT7_Mn7@1025_d N_OUT6_Mn7@1025_g N_VSS_Mn7@1025_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1024 N_OUT7_Mn7@1024_d N_OUT6_Mn7@1024_g N_VSS_Mn7@1024_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1025 N_OUT7_Mp7@1025_d N_OUT6_Mp7@1025_g N_VDD_Mp7@1025_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1024 N_OUT7_Mp7@1024_d N_OUT6_Mp7@1024_g N_VDD_Mp7@1024_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1023 N_OUT7_Mn7@1023_d N_OUT6_Mn7@1023_g N_VSS_Mn7@1023_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1022 N_OUT7_Mn7@1022_d N_OUT6_Mn7@1022_g N_VSS_Mn7@1022_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1023 N_OUT7_Mp7@1023_d N_OUT6_Mp7@1023_g N_VDD_Mp7@1023_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1022 N_OUT7_Mp7@1022_d N_OUT6_Mp7@1022_g N_VDD_Mp7@1022_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1021 N_OUT7_Mn7@1021_d N_OUT6_Mn7@1021_g N_VSS_Mn7@1021_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1020 N_OUT7_Mn7@1020_d N_OUT6_Mn7@1020_g N_VSS_Mn7@1020_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1021 N_OUT7_Mp7@1021_d N_OUT6_Mp7@1021_g N_VDD_Mp7@1021_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1020 N_OUT7_Mp7@1020_d N_OUT6_Mp7@1020_g N_VDD_Mp7@1020_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1019 N_OUT7_Mn7@1019_d N_OUT6_Mn7@1019_g N_VSS_Mn7@1019_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1018 N_OUT7_Mn7@1018_d N_OUT6_Mn7@1018_g N_VSS_Mn7@1018_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1019 N_OUT7_Mp7@1019_d N_OUT6_Mp7@1019_g N_VDD_Mp7@1019_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1018 N_OUT7_Mp7@1018_d N_OUT6_Mp7@1018_g N_VDD_Mp7@1018_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1017 N_OUT7_Mn7@1017_d N_OUT6_Mn7@1017_g N_VSS_Mn7@1017_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1016 N_OUT7_Mn7@1016_d N_OUT6_Mn7@1016_g N_VSS_Mn7@1016_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1017 N_OUT7_Mp7@1017_d N_OUT6_Mp7@1017_g N_VDD_Mp7@1017_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1016 N_OUT7_Mp7@1016_d N_OUT6_Mp7@1016_g N_VDD_Mp7@1016_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1015 N_OUT7_Mn7@1015_d N_OUT6_Mn7@1015_g N_VSS_Mn7@1015_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1014 N_OUT7_Mn7@1014_d N_OUT6_Mn7@1014_g N_VSS_Mn7@1014_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1015 N_OUT7_Mp7@1015_d N_OUT6_Mp7@1015_g N_VDD_Mp7@1015_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1014 N_OUT7_Mp7@1014_d N_OUT6_Mp7@1014_g N_VDD_Mp7@1014_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1013 N_OUT7_Mn7@1013_d N_OUT6_Mn7@1013_g N_VSS_Mn7@1013_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1012 N_OUT7_Mn7@1012_d N_OUT6_Mn7@1012_g N_VSS_Mn7@1012_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1013 N_OUT7_Mp7@1013_d N_OUT6_Mp7@1013_g N_VDD_Mp7@1013_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1012 N_OUT7_Mp7@1012_d N_OUT6_Mp7@1012_g N_VDD_Mp7@1012_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1011 N_OUT7_Mn7@1011_d N_OUT6_Mn7@1011_g N_VSS_Mn7@1011_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1010 N_OUT7_Mn7@1010_d N_OUT6_Mn7@1010_g N_VSS_Mn7@1010_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1011 N_OUT7_Mp7@1011_d N_OUT6_Mp7@1011_g N_VDD_Mp7@1011_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1010 N_OUT7_Mp7@1010_d N_OUT6_Mp7@1010_g N_VDD_Mp7@1010_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1009 N_OUT7_Mn7@1009_d N_OUT6_Mn7@1009_g N_VSS_Mn7@1009_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1008 N_OUT7_Mn7@1008_d N_OUT6_Mn7@1008_g N_VSS_Mn7@1008_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1009 N_OUT7_Mp7@1009_d N_OUT6_Mp7@1009_g N_VDD_Mp7@1009_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1008 N_OUT7_Mp7@1008_d N_OUT6_Mp7@1008_g N_VDD_Mp7@1008_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1007 N_OUT7_Mn7@1007_d N_OUT6_Mn7@1007_g N_VSS_Mn7@1007_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1006 N_OUT7_Mn7@1006_d N_OUT6_Mn7@1006_g N_VSS_Mn7@1006_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1007 N_OUT7_Mp7@1007_d N_OUT6_Mp7@1007_g N_VDD_Mp7@1007_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1006 N_OUT7_Mp7@1006_d N_OUT6_Mp7@1006_g N_VDD_Mp7@1006_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1005 N_OUT7_Mn7@1005_d N_OUT6_Mn7@1005_g N_VSS_Mn7@1005_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1004 N_OUT7_Mn7@1004_d N_OUT6_Mn7@1004_g N_VSS_Mn7@1004_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1005 N_OUT7_Mp7@1005_d N_OUT6_Mp7@1005_g N_VDD_Mp7@1005_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1004 N_OUT7_Mp7@1004_d N_OUT6_Mp7@1004_g N_VDD_Mp7@1004_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1003 N_OUT7_Mn7@1003_d N_OUT6_Mn7@1003_g N_VSS_Mn7@1003_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1002 N_OUT7_Mn7@1002_d N_OUT6_Mn7@1002_g N_VSS_Mn7@1002_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1003 N_OUT7_Mp7@1003_d N_OUT6_Mp7@1003_g N_VDD_Mp7@1003_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1002 N_OUT7_Mp7@1002_d N_OUT6_Mp7@1002_g N_VDD_Mp7@1002_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@1001 N_OUT7_Mn7@1001_d N_OUT6_Mn7@1001_g N_VSS_Mn7@1001_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@1000 N_OUT7_Mn7@1000_d N_OUT6_Mn7@1000_g N_VSS_Mn7@1000_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@1001 N_OUT7_Mp7@1001_d N_OUT6_Mp7@1001_g N_VDD_Mp7@1001_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@1000 N_OUT7_Mp7@1000_d N_OUT6_Mp7@1000_g N_VDD_Mp7@1000_s N_VDD_Mp7@1159_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@999 N_OUT7_Mn7@999_d N_OUT6_Mn7@999_g N_VSS_Mn7@999_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@998 N_OUT7_Mn7@998_d N_OUT6_Mn7@998_g N_VSS_Mn7@998_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@999 N_OUT7_Mp7@999_d N_OUT6_Mp7@999_g N_VDD_Mp7@999_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@998 N_OUT7_Mp7@998_d N_OUT6_Mp7@998_g N_VDD_Mp7@998_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@997 N_OUT7_Mn7@997_d N_OUT6_Mn7@997_g N_VSS_Mn7@997_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@996 N_OUT7_Mn7@996_d N_OUT6_Mn7@996_g N_VSS_Mn7@996_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@997 N_OUT7_Mp7@997_d N_OUT6_Mp7@997_g N_VDD_Mp7@997_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@996 N_OUT7_Mp7@996_d N_OUT6_Mp7@996_g N_VDD_Mp7@996_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@995 N_OUT7_Mn7@995_d N_OUT6_Mn7@995_g N_VSS_Mn7@995_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@994 N_OUT7_Mn7@994_d N_OUT6_Mn7@994_g N_VSS_Mn7@994_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@995 N_OUT7_Mp7@995_d N_OUT6_Mp7@995_g N_VDD_Mp7@995_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@994 N_OUT7_Mp7@994_d N_OUT6_Mp7@994_g N_VDD_Mp7@994_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@993 N_OUT7_Mn7@993_d N_OUT6_Mn7@993_g N_VSS_Mn7@993_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@992 N_OUT7_Mn7@992_d N_OUT6_Mn7@992_g N_VSS_Mn7@992_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@993 N_OUT7_Mp7@993_d N_OUT6_Mp7@993_g N_VDD_Mp7@993_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@992 N_OUT7_Mp7@992_d N_OUT6_Mp7@992_g N_VDD_Mp7@992_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@991 N_OUT7_Mn7@991_d N_OUT6_Mn7@991_g N_VSS_Mn7@991_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@990 N_OUT7_Mn7@990_d N_OUT6_Mn7@990_g N_VSS_Mn7@990_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@991 N_OUT7_Mp7@991_d N_OUT6_Mp7@991_g N_VDD_Mp7@991_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@990 N_OUT7_Mp7@990_d N_OUT6_Mp7@990_g N_VDD_Mp7@990_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@989 N_OUT7_Mn7@989_d N_OUT6_Mn7@989_g N_VSS_Mn7@989_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@988 N_OUT7_Mn7@988_d N_OUT6_Mn7@988_g N_VSS_Mn7@988_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@989 N_OUT7_Mp7@989_d N_OUT6_Mp7@989_g N_VDD_Mp7@989_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@988 N_OUT7_Mp7@988_d N_OUT6_Mp7@988_g N_VDD_Mp7@988_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@987 N_OUT7_Mn7@987_d N_OUT6_Mn7@987_g N_VSS_Mn7@987_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@986 N_OUT7_Mn7@986_d N_OUT6_Mn7@986_g N_VSS_Mn7@986_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@987 N_OUT7_Mp7@987_d N_OUT6_Mp7@987_g N_VDD_Mp7@987_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@986 N_OUT7_Mp7@986_d N_OUT6_Mp7@986_g N_VDD_Mp7@986_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@985 N_OUT7_Mn7@985_d N_OUT6_Mn7@985_g N_VSS_Mn7@985_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@984 N_OUT7_Mn7@984_d N_OUT6_Mn7@984_g N_VSS_Mn7@984_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@985 N_OUT7_Mp7@985_d N_OUT6_Mp7@985_g N_VDD_Mp7@985_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@984 N_OUT7_Mp7@984_d N_OUT6_Mp7@984_g N_VDD_Mp7@984_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@983 N_OUT7_Mn7@983_d N_OUT6_Mn7@983_g N_VSS_Mn7@983_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@982 N_OUT7_Mn7@982_d N_OUT6_Mn7@982_g N_VSS_Mn7@982_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@983 N_OUT7_Mp7@983_d N_OUT6_Mp7@983_g N_VDD_Mp7@983_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@982 N_OUT7_Mp7@982_d N_OUT6_Mp7@982_g N_VDD_Mp7@982_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@981 N_OUT7_Mn7@981_d N_OUT6_Mn7@981_g N_VSS_Mn7@981_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@980 N_OUT7_Mn7@980_d N_OUT6_Mn7@980_g N_VSS_Mn7@980_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@981 N_OUT7_Mp7@981_d N_OUT6_Mp7@981_g N_VDD_Mp7@981_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@980 N_OUT7_Mp7@980_d N_OUT6_Mp7@980_g N_VDD_Mp7@980_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@979 N_OUT7_Mn7@979_d N_OUT6_Mn7@979_g N_VSS_Mn7@979_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@978 N_OUT7_Mn7@978_d N_OUT6_Mn7@978_g N_VSS_Mn7@978_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@979 N_OUT7_Mp7@979_d N_OUT6_Mp7@979_g N_VDD_Mp7@979_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@978 N_OUT7_Mp7@978_d N_OUT6_Mp7@978_g N_VDD_Mp7@978_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@977 N_OUT7_Mn7@977_d N_OUT6_Mn7@977_g N_VSS_Mn7@977_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@976 N_OUT7_Mn7@976_d N_OUT6_Mn7@976_g N_VSS_Mn7@976_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@977 N_OUT7_Mp7@977_d N_OUT6_Mp7@977_g N_VDD_Mp7@977_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@976 N_OUT7_Mp7@976_d N_OUT6_Mp7@976_g N_VDD_Mp7@976_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@975 N_OUT7_Mn7@975_d N_OUT6_Mn7@975_g N_VSS_Mn7@975_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@974 N_OUT7_Mn7@974_d N_OUT6_Mn7@974_g N_VSS_Mn7@974_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@975 N_OUT7_Mp7@975_d N_OUT6_Mp7@975_g N_VDD_Mp7@975_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@974 N_OUT7_Mp7@974_d N_OUT6_Mp7@974_g N_VDD_Mp7@974_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@973 N_OUT7_Mn7@973_d N_OUT6_Mn7@973_g N_VSS_Mn7@973_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@972 N_OUT7_Mn7@972_d N_OUT6_Mn7@972_g N_VSS_Mn7@972_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@973 N_OUT7_Mp7@973_d N_OUT6_Mp7@973_g N_VDD_Mp7@973_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@972 N_OUT7_Mp7@972_d N_OUT6_Mp7@972_g N_VDD_Mp7@972_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@971 N_OUT7_Mn7@971_d N_OUT6_Mn7@971_g N_VSS_Mn7@971_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@970 N_OUT7_Mn7@970_d N_OUT6_Mn7@970_g N_VSS_Mn7@970_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@971 N_OUT7_Mp7@971_d N_OUT6_Mp7@971_g N_VDD_Mp7@971_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@970 N_OUT7_Mp7@970_d N_OUT6_Mp7@970_g N_VDD_Mp7@970_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@969 N_OUT7_Mn7@969_d N_OUT6_Mn7@969_g N_VSS_Mn7@969_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@968 N_OUT7_Mn7@968_d N_OUT6_Mn7@968_g N_VSS_Mn7@968_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@969 N_OUT7_Mp7@969_d N_OUT6_Mp7@969_g N_VDD_Mp7@969_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@968 N_OUT7_Mp7@968_d N_OUT6_Mp7@968_g N_VDD_Mp7@968_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@967 N_OUT7_Mn7@967_d N_OUT6_Mn7@967_g N_VSS_Mn7@967_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@966 N_OUT7_Mn7@966_d N_OUT6_Mn7@966_g N_VSS_Mn7@966_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@967 N_OUT7_Mp7@967_d N_OUT6_Mp7@967_g N_VDD_Mp7@967_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@966 N_OUT7_Mp7@966_d N_OUT6_Mp7@966_g N_VDD_Mp7@966_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@965 N_OUT7_Mn7@965_d N_OUT6_Mn7@965_g N_VSS_Mn7@965_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@964 N_OUT7_Mn7@964_d N_OUT6_Mn7@964_g N_VSS_Mn7@964_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@965 N_OUT7_Mp7@965_d N_OUT6_Mp7@965_g N_VDD_Mp7@965_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@964 N_OUT7_Mp7@964_d N_OUT6_Mp7@964_g N_VDD_Mp7@964_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@963 N_OUT7_Mn7@963_d N_OUT6_Mn7@963_g N_VSS_Mn7@963_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@962 N_OUT7_Mn7@962_d N_OUT6_Mn7@962_g N_VSS_Mn7@962_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@963 N_OUT7_Mp7@963_d N_OUT6_Mp7@963_g N_VDD_Mp7@963_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@962 N_OUT7_Mp7@962_d N_OUT6_Mp7@962_g N_VDD_Mp7@962_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@961 N_OUT7_Mn7@961_d N_OUT6_Mn7@961_g N_VSS_Mn7@961_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@960 N_OUT7_Mn7@960_d N_OUT6_Mn7@960_g N_VSS_Mn7@960_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@961 N_OUT7_Mp7@961_d N_OUT6_Mp7@961_g N_VDD_Mp7@961_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@960 N_OUT7_Mp7@960_d N_OUT6_Mp7@960_g N_VDD_Mp7@960_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@959 N_OUT7_Mn7@959_d N_OUT6_Mn7@959_g N_VSS_Mn7@959_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@958 N_OUT7_Mn7@958_d N_OUT6_Mn7@958_g N_VSS_Mn7@958_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@959 N_OUT7_Mp7@959_d N_OUT6_Mp7@959_g N_VDD_Mp7@959_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@958 N_OUT7_Mp7@958_d N_OUT6_Mp7@958_g N_VDD_Mp7@958_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@957 N_OUT7_Mn7@957_d N_OUT6_Mn7@957_g N_VSS_Mn7@957_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@956 N_OUT7_Mn7@956_d N_OUT6_Mn7@956_g N_VSS_Mn7@956_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@957 N_OUT7_Mp7@957_d N_OUT6_Mp7@957_g N_VDD_Mp7@957_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@956 N_OUT7_Mp7@956_d N_OUT6_Mp7@956_g N_VDD_Mp7@956_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@955 N_OUT7_Mn7@955_d N_OUT6_Mn7@955_g N_VSS_Mn7@955_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@954 N_OUT7_Mn7@954_d N_OUT6_Mn7@954_g N_VSS_Mn7@954_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@955 N_OUT7_Mp7@955_d N_OUT6_Mp7@955_g N_VDD_Mp7@955_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@954 N_OUT7_Mp7@954_d N_OUT6_Mp7@954_g N_VDD_Mp7@954_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@953 N_OUT7_Mn7@953_d N_OUT6_Mn7@953_g N_VSS_Mn7@953_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@952 N_OUT7_Mn7@952_d N_OUT6_Mn7@952_g N_VSS_Mn7@952_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@953 N_OUT7_Mp7@953_d N_OUT6_Mp7@953_g N_VDD_Mp7@953_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@952 N_OUT7_Mp7@952_d N_OUT6_Mp7@952_g N_VDD_Mp7@952_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@951 N_OUT7_Mn7@951_d N_OUT6_Mn7@951_g N_VSS_Mn7@951_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@950 N_OUT7_Mn7@950_d N_OUT6_Mn7@950_g N_VSS_Mn7@950_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@951 N_OUT7_Mp7@951_d N_OUT6_Mp7@951_g N_VDD_Mp7@951_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@950 N_OUT7_Mp7@950_d N_OUT6_Mp7@950_g N_VDD_Mp7@950_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@949 N_OUT7_Mn7@949_d N_OUT6_Mn7@949_g N_VSS_Mn7@949_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@948 N_OUT7_Mn7@948_d N_OUT6_Mn7@948_g N_VSS_Mn7@948_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@949 N_OUT7_Mp7@949_d N_OUT6_Mp7@949_g N_VDD_Mp7@949_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@948 N_OUT7_Mp7@948_d N_OUT6_Mp7@948_g N_VDD_Mp7@948_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@947 N_OUT7_Mn7@947_d N_OUT6_Mn7@947_g N_VSS_Mn7@947_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@946 N_OUT7_Mn7@946_d N_OUT6_Mn7@946_g N_VSS_Mn7@946_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@947 N_OUT7_Mp7@947_d N_OUT6_Mp7@947_g N_VDD_Mp7@947_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@946 N_OUT7_Mp7@946_d N_OUT6_Mp7@946_g N_VDD_Mp7@946_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@945 N_OUT7_Mn7@945_d N_OUT6_Mn7@945_g N_VSS_Mn7@945_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@944 N_OUT7_Mn7@944_d N_OUT6_Mn7@944_g N_VSS_Mn7@944_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@945 N_OUT7_Mp7@945_d N_OUT6_Mp7@945_g N_VDD_Mp7@945_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@944 N_OUT7_Mp7@944_d N_OUT6_Mp7@944_g N_VDD_Mp7@944_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@943 N_OUT7_Mn7@943_d N_OUT6_Mn7@943_g N_VSS_Mn7@943_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@942 N_OUT7_Mn7@942_d N_OUT6_Mn7@942_g N_VSS_Mn7@942_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@943 N_OUT7_Mp7@943_d N_OUT6_Mp7@943_g N_VDD_Mp7@943_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@942 N_OUT7_Mp7@942_d N_OUT6_Mp7@942_g N_VDD_Mp7@942_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@941 N_OUT7_Mn7@941_d N_OUT6_Mn7@941_g N_VSS_Mn7@941_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@940 N_OUT7_Mn7@940_d N_OUT6_Mn7@940_g N_VSS_Mn7@940_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@941 N_OUT7_Mp7@941_d N_OUT6_Mp7@941_g N_VDD_Mp7@941_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@940 N_OUT7_Mp7@940_d N_OUT6_Mp7@940_g N_VDD_Mp7@940_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@939 N_OUT7_Mn7@939_d N_OUT6_Mn7@939_g N_VSS_Mn7@939_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@938 N_OUT7_Mn7@938_d N_OUT6_Mn7@938_g N_VSS_Mn7@938_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@939 N_OUT7_Mp7@939_d N_OUT6_Mp7@939_g N_VDD_Mp7@939_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@938 N_OUT7_Mp7@938_d N_OUT6_Mp7@938_g N_VDD_Mp7@938_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@937 N_OUT7_Mn7@937_d N_OUT6_Mn7@937_g N_VSS_Mn7@937_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@936 N_OUT7_Mn7@936_d N_OUT6_Mn7@936_g N_VSS_Mn7@936_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@937 N_OUT7_Mp7@937_d N_OUT6_Mp7@937_g N_VDD_Mp7@937_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@936 N_OUT7_Mp7@936_d N_OUT6_Mp7@936_g N_VDD_Mp7@936_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@935 N_OUT7_Mn7@935_d N_OUT6_Mn7@935_g N_VSS_Mn7@935_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@934 N_OUT7_Mn7@934_d N_OUT6_Mn7@934_g N_VSS_Mn7@934_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@935 N_OUT7_Mp7@935_d N_OUT6_Mp7@935_g N_VDD_Mp7@935_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@934 N_OUT7_Mp7@934_d N_OUT6_Mp7@934_g N_VDD_Mp7@934_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@933 N_OUT7_Mn7@933_d N_OUT6_Mn7@933_g N_VSS_Mn7@933_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@932 N_OUT7_Mn7@932_d N_OUT6_Mn7@932_g N_VSS_Mn7@932_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@933 N_OUT7_Mp7@933_d N_OUT6_Mp7@933_g N_VDD_Mp7@933_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@932 N_OUT7_Mp7@932_d N_OUT6_Mp7@932_g N_VDD_Mp7@932_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@931 N_OUT7_Mn7@931_d N_OUT6_Mn7@931_g N_VSS_Mn7@931_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@930 N_OUT7_Mn7@930_d N_OUT6_Mn7@930_g N_VSS_Mn7@930_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@931 N_OUT7_Mp7@931_d N_OUT6_Mp7@931_g N_VDD_Mp7@931_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@930 N_OUT7_Mp7@930_d N_OUT6_Mp7@930_g N_VDD_Mp7@930_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@929 N_OUT7_Mn7@929_d N_OUT6_Mn7@929_g N_VSS_Mn7@929_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@928 N_OUT7_Mn7@928_d N_OUT6_Mn7@928_g N_VSS_Mn7@928_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@929 N_OUT7_Mp7@929_d N_OUT6_Mp7@929_g N_VDD_Mp7@929_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@928 N_OUT7_Mp7@928_d N_OUT6_Mp7@928_g N_VDD_Mp7@928_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@927 N_OUT7_Mn7@927_d N_OUT6_Mn7@927_g N_VSS_Mn7@927_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@926 N_OUT7_Mn7@926_d N_OUT6_Mn7@926_g N_VSS_Mn7@926_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@927 N_OUT7_Mp7@927_d N_OUT6_Mp7@927_g N_VDD_Mp7@927_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@926 N_OUT7_Mp7@926_d N_OUT6_Mp7@926_g N_VDD_Mp7@926_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@925 N_OUT7_Mn7@925_d N_OUT6_Mn7@925_g N_VSS_Mn7@925_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@924 N_OUT7_Mn7@924_d N_OUT6_Mn7@924_g N_VSS_Mn7@924_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@925 N_OUT7_Mp7@925_d N_OUT6_Mp7@925_g N_VDD_Mp7@925_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@924 N_OUT7_Mp7@924_d N_OUT6_Mp7@924_g N_VDD_Mp7@924_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@923 N_OUT7_Mn7@923_d N_OUT6_Mn7@923_g N_VSS_Mn7@923_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@922 N_OUT7_Mn7@922_d N_OUT6_Mn7@922_g N_VSS_Mn7@922_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@923 N_OUT7_Mp7@923_d N_OUT6_Mp7@923_g N_VDD_Mp7@923_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@922 N_OUT7_Mp7@922_d N_OUT6_Mp7@922_g N_VDD_Mp7@922_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@921 N_OUT7_Mn7@921_d N_OUT6_Mn7@921_g N_VSS_Mn7@921_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@920 N_OUT7_Mn7@920_d N_OUT6_Mn7@920_g N_VSS_Mn7@920_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@921 N_OUT7_Mp7@921_d N_OUT6_Mp7@921_g N_VDD_Mp7@921_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@920 N_OUT7_Mp7@920_d N_OUT6_Mp7@920_g N_VDD_Mp7@920_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@919 N_OUT7_Mn7@919_d N_OUT6_Mn7@919_g N_VSS_Mn7@919_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@918 N_OUT7_Mn7@918_d N_OUT6_Mn7@918_g N_VSS_Mn7@918_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@919 N_OUT7_Mp7@919_d N_OUT6_Mp7@919_g N_VDD_Mp7@919_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@918 N_OUT7_Mp7@918_d N_OUT6_Mp7@918_g N_VDD_Mp7@918_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@917 N_OUT7_Mn7@917_d N_OUT6_Mn7@917_g N_VSS_Mn7@917_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@916 N_OUT7_Mn7@916_d N_OUT6_Mn7@916_g N_VSS_Mn7@916_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@917 N_OUT7_Mp7@917_d N_OUT6_Mp7@917_g N_VDD_Mp7@917_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@916 N_OUT7_Mp7@916_d N_OUT6_Mp7@916_g N_VDD_Mp7@916_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@915 N_OUT7_Mn7@915_d N_OUT6_Mn7@915_g N_VSS_Mn7@915_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@914 N_OUT7_Mn7@914_d N_OUT6_Mn7@914_g N_VSS_Mn7@914_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@915 N_OUT7_Mp7@915_d N_OUT6_Mp7@915_g N_VDD_Mp7@915_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@914 N_OUT7_Mp7@914_d N_OUT6_Mp7@914_g N_VDD_Mp7@914_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@913 N_OUT7_Mn7@913_d N_OUT6_Mn7@913_g N_VSS_Mn7@913_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@912 N_OUT7_Mn7@912_d N_OUT6_Mn7@912_g N_VSS_Mn7@912_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@913 N_OUT7_Mp7@913_d N_OUT6_Mp7@913_g N_VDD_Mp7@913_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@912 N_OUT7_Mp7@912_d N_OUT6_Mp7@912_g N_VDD_Mp7@912_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@911 N_OUT7_Mn7@911_d N_OUT6_Mn7@911_g N_VSS_Mn7@911_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@910 N_OUT7_Mn7@910_d N_OUT6_Mn7@910_g N_VSS_Mn7@910_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@911 N_OUT7_Mp7@911_d N_OUT6_Mp7@911_g N_VDD_Mp7@911_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@910 N_OUT7_Mp7@910_d N_OUT6_Mp7@910_g N_VDD_Mp7@910_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@909 N_OUT7_Mn7@909_d N_OUT6_Mn7@909_g N_VSS_Mn7@909_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@908 N_OUT7_Mn7@908_d N_OUT6_Mn7@908_g N_VSS_Mn7@908_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@909 N_OUT7_Mp7@909_d N_OUT6_Mp7@909_g N_VDD_Mp7@909_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@908 N_OUT7_Mp7@908_d N_OUT6_Mp7@908_g N_VDD_Mp7@908_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@907 N_OUT7_Mn7@907_d N_OUT6_Mn7@907_g N_VSS_Mn7@907_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@906 N_OUT7_Mn7@906_d N_OUT6_Mn7@906_g N_VSS_Mn7@906_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@907 N_OUT7_Mp7@907_d N_OUT6_Mp7@907_g N_VDD_Mp7@907_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@906 N_OUT7_Mp7@906_d N_OUT6_Mp7@906_g N_VDD_Mp7@906_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@905 N_OUT7_Mn7@905_d N_OUT6_Mn7@905_g N_VSS_Mn7@905_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@904 N_OUT7_Mn7@904_d N_OUT6_Mn7@904_g N_VSS_Mn7@904_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@905 N_OUT7_Mp7@905_d N_OUT6_Mp7@905_g N_VDD_Mp7@905_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@904 N_OUT7_Mp7@904_d N_OUT6_Mp7@904_g N_VDD_Mp7@904_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@903 N_OUT7_Mn7@903_d N_OUT6_Mn7@903_g N_VSS_Mn7@903_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@902 N_OUT7_Mn7@902_d N_OUT6_Mn7@902_g N_VSS_Mn7@902_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@903 N_OUT7_Mp7@903_d N_OUT6_Mp7@903_g N_VDD_Mp7@903_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@902 N_OUT7_Mp7@902_d N_OUT6_Mp7@902_g N_VDD_Mp7@902_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@901 N_OUT7_Mn7@901_d N_OUT6_Mn7@901_g N_VSS_Mn7@901_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@900 N_OUT7_Mn7@900_d N_OUT6_Mn7@900_g N_VSS_Mn7@900_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@901 N_OUT7_Mp7@901_d N_OUT6_Mp7@901_g N_VDD_Mp7@901_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@900 N_OUT7_Mp7@900_d N_OUT6_Mp7@900_g N_VDD_Mp7@900_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@899 N_OUT7_Mn7@899_d N_OUT6_Mn7@899_g N_VSS_Mn7@899_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@898 N_OUT7_Mn7@898_d N_OUT6_Mn7@898_g N_VSS_Mn7@898_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@899 N_OUT7_Mp7@899_d N_OUT6_Mp7@899_g N_VDD_Mp7@899_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@898 N_OUT7_Mp7@898_d N_OUT6_Mp7@898_g N_VDD_Mp7@898_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@897 N_OUT7_Mn7@897_d N_OUT6_Mn7@897_g N_VSS_Mn7@897_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@896 N_OUT7_Mn7@896_d N_OUT6_Mn7@896_g N_VSS_Mn7@896_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@897 N_OUT7_Mp7@897_d N_OUT6_Mp7@897_g N_VDD_Mp7@897_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@896 N_OUT7_Mp7@896_d N_OUT6_Mp7@896_g N_VDD_Mp7@896_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@895 N_OUT7_Mn7@895_d N_OUT6_Mn7@895_g N_VSS_Mn7@895_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@894 N_OUT7_Mn7@894_d N_OUT6_Mn7@894_g N_VSS_Mn7@894_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@895 N_OUT7_Mp7@895_d N_OUT6_Mp7@895_g N_VDD_Mp7@895_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@894 N_OUT7_Mp7@894_d N_OUT6_Mp7@894_g N_VDD_Mp7@894_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@893 N_OUT7_Mn7@893_d N_OUT6_Mn7@893_g N_VSS_Mn7@893_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@892 N_OUT7_Mn7@892_d N_OUT6_Mn7@892_g N_VSS_Mn7@892_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@893 N_OUT7_Mp7@893_d N_OUT6_Mp7@893_g N_VDD_Mp7@893_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@892 N_OUT7_Mp7@892_d N_OUT6_Mp7@892_g N_VDD_Mp7@892_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@891 N_OUT7_Mn7@891_d N_OUT6_Mn7@891_g N_VSS_Mn7@891_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@890 N_OUT7_Mn7@890_d N_OUT6_Mn7@890_g N_VSS_Mn7@890_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@891 N_OUT7_Mp7@891_d N_OUT6_Mp7@891_g N_VDD_Mp7@891_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@890 N_OUT7_Mp7@890_d N_OUT6_Mp7@890_g N_VDD_Mp7@890_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@889 N_OUT7_Mn7@889_d N_OUT6_Mn7@889_g N_VSS_Mn7@889_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@888 N_OUT7_Mn7@888_d N_OUT6_Mn7@888_g N_VSS_Mn7@888_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@889 N_OUT7_Mp7@889_d N_OUT6_Mp7@889_g N_VDD_Mp7@889_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@888 N_OUT7_Mp7@888_d N_OUT6_Mp7@888_g N_VDD_Mp7@888_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@887 N_OUT7_Mn7@887_d N_OUT6_Mn7@887_g N_VSS_Mn7@887_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@886 N_OUT7_Mn7@886_d N_OUT6_Mn7@886_g N_VSS_Mn7@886_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@887 N_OUT7_Mp7@887_d N_OUT6_Mp7@887_g N_VDD_Mp7@887_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@886 N_OUT7_Mp7@886_d N_OUT6_Mp7@886_g N_VDD_Mp7@886_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@885 N_OUT7_Mn7@885_d N_OUT6_Mn7@885_g N_VSS_Mn7@885_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@884 N_OUT7_Mn7@884_d N_OUT6_Mn7@884_g N_VSS_Mn7@884_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@885 N_OUT7_Mp7@885_d N_OUT6_Mp7@885_g N_VDD_Mp7@885_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@884 N_OUT7_Mp7@884_d N_OUT6_Mp7@884_g N_VDD_Mp7@884_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@883 N_OUT7_Mn7@883_d N_OUT6_Mn7@883_g N_VSS_Mn7@883_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@882 N_OUT7_Mn7@882_d N_OUT6_Mn7@882_g N_VSS_Mn7@882_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@883 N_OUT7_Mp7@883_d N_OUT6_Mp7@883_g N_VDD_Mp7@883_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@882 N_OUT7_Mp7@882_d N_OUT6_Mp7@882_g N_VDD_Mp7@882_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@881 N_OUT7_Mn7@881_d N_OUT6_Mn7@881_g N_VSS_Mn7@881_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@880 N_OUT7_Mn7@880_d N_OUT6_Mn7@880_g N_VSS_Mn7@880_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@881 N_OUT7_Mp7@881_d N_OUT6_Mp7@881_g N_VDD_Mp7@881_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@880 N_OUT7_Mp7@880_d N_OUT6_Mp7@880_g N_VDD_Mp7@880_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@879 N_OUT7_Mn7@879_d N_OUT6_Mn7@879_g N_VSS_Mn7@879_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@878 N_OUT7_Mn7@878_d N_OUT6_Mn7@878_g N_VSS_Mn7@878_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@879 N_OUT7_Mp7@879_d N_OUT6_Mp7@879_g N_VDD_Mp7@879_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@878 N_OUT7_Mp7@878_d N_OUT6_Mp7@878_g N_VDD_Mp7@878_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@877 N_OUT7_Mn7@877_d N_OUT6_Mn7@877_g N_VSS_Mn7@877_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@876 N_OUT7_Mn7@876_d N_OUT6_Mn7@876_g N_VSS_Mn7@876_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@877 N_OUT7_Mp7@877_d N_OUT6_Mp7@877_g N_VDD_Mp7@877_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@876 N_OUT7_Mp7@876_d N_OUT6_Mp7@876_g N_VDD_Mp7@876_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@875 N_OUT7_Mn7@875_d N_OUT6_Mn7@875_g N_VSS_Mn7@875_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@874 N_OUT7_Mn7@874_d N_OUT6_Mn7@874_g N_VSS_Mn7@874_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@875 N_OUT7_Mp7@875_d N_OUT6_Mp7@875_g N_VDD_Mp7@875_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@874 N_OUT7_Mp7@874_d N_OUT6_Mp7@874_g N_VDD_Mp7@874_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@873 N_OUT7_Mn7@873_d N_OUT6_Mn7@873_g N_VSS_Mn7@873_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@872 N_OUT7_Mn7@872_d N_OUT6_Mn7@872_g N_VSS_Mn7@872_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@873 N_OUT7_Mp7@873_d N_OUT6_Mp7@873_g N_VDD_Mp7@873_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@872 N_OUT7_Mp7@872_d N_OUT6_Mp7@872_g N_VDD_Mp7@872_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@871 N_OUT7_Mn7@871_d N_OUT6_Mn7@871_g N_VSS_Mn7@871_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@870 N_OUT7_Mn7@870_d N_OUT6_Mn7@870_g N_VSS_Mn7@870_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@871 N_OUT7_Mp7@871_d N_OUT6_Mp7@871_g N_VDD_Mp7@871_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@870 N_OUT7_Mp7@870_d N_OUT6_Mp7@870_g N_VDD_Mp7@870_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@869 N_OUT7_Mn7@869_d N_OUT6_Mn7@869_g N_VSS_Mn7@869_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@868 N_OUT7_Mn7@868_d N_OUT6_Mn7@868_g N_VSS_Mn7@868_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@869 N_OUT7_Mp7@869_d N_OUT6_Mp7@869_g N_VDD_Mp7@869_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@868 N_OUT7_Mp7@868_d N_OUT6_Mp7@868_g N_VDD_Mp7@868_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@867 N_OUT7_Mn7@867_d N_OUT6_Mn7@867_g N_VSS_Mn7@867_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@866 N_OUT7_Mn7@866_d N_OUT6_Mn7@866_g N_VSS_Mn7@866_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@867 N_OUT7_Mp7@867_d N_OUT6_Mp7@867_g N_VDD_Mp7@867_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@866 N_OUT7_Mp7@866_d N_OUT6_Mp7@866_g N_VDD_Mp7@866_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@865 N_OUT7_Mn7@865_d N_OUT6_Mn7@865_g N_VSS_Mn7@865_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@864 N_OUT7_Mn7@864_d N_OUT6_Mn7@864_g N_VSS_Mn7@864_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@865 N_OUT7_Mp7@865_d N_OUT6_Mp7@865_g N_VDD_Mp7@865_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@864 N_OUT7_Mp7@864_d N_OUT6_Mp7@864_g N_VDD_Mp7@864_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@863 N_OUT7_Mn7@863_d N_OUT6_Mn7@863_g N_VSS_Mn7@863_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@862 N_OUT7_Mn7@862_d N_OUT6_Mn7@862_g N_VSS_Mn7@862_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@863 N_OUT7_Mp7@863_d N_OUT6_Mp7@863_g N_VDD_Mp7@863_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@862 N_OUT7_Mp7@862_d N_OUT6_Mp7@862_g N_VDD_Mp7@862_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@861 N_OUT7_Mn7@861_d N_OUT6_Mn7@861_g N_VSS_Mn7@861_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@860 N_OUT7_Mn7@860_d N_OUT6_Mn7@860_g N_VSS_Mn7@860_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@861 N_OUT7_Mp7@861_d N_OUT6_Mp7@861_g N_VDD_Mp7@861_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@860 N_OUT7_Mp7@860_d N_OUT6_Mp7@860_g N_VDD_Mp7@860_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@859 N_OUT7_Mn7@859_d N_OUT6_Mn7@859_g N_VSS_Mn7@859_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@858 N_OUT7_Mn7@858_d N_OUT6_Mn7@858_g N_VSS_Mn7@858_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@859 N_OUT7_Mp7@859_d N_OUT6_Mp7@859_g N_VDD_Mp7@859_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@858 N_OUT7_Mp7@858_d N_OUT6_Mp7@858_g N_VDD_Mp7@858_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@857 N_OUT7_Mn7@857_d N_OUT6_Mn7@857_g N_VSS_Mn7@857_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@856 N_OUT7_Mn7@856_d N_OUT6_Mn7@856_g N_VSS_Mn7@856_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@857 N_OUT7_Mp7@857_d N_OUT6_Mp7@857_g N_VDD_Mp7@857_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@856 N_OUT7_Mp7@856_d N_OUT6_Mp7@856_g N_VDD_Mp7@856_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@855 N_OUT7_Mn7@855_d N_OUT6_Mn7@855_g N_VSS_Mn7@855_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@854 N_OUT7_Mn7@854_d N_OUT6_Mn7@854_g N_VSS_Mn7@854_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@855 N_OUT7_Mp7@855_d N_OUT6_Mp7@855_g N_VDD_Mp7@855_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@854 N_OUT7_Mp7@854_d N_OUT6_Mp7@854_g N_VDD_Mp7@854_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@853 N_OUT7_Mn7@853_d N_OUT6_Mn7@853_g N_VSS_Mn7@853_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@852 N_OUT7_Mn7@852_d N_OUT6_Mn7@852_g N_VSS_Mn7@852_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@853 N_OUT7_Mp7@853_d N_OUT6_Mp7@853_g N_VDD_Mp7@853_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@852 N_OUT7_Mp7@852_d N_OUT6_Mp7@852_g N_VDD_Mp7@852_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@851 N_OUT7_Mn7@851_d N_OUT6_Mn7@851_g N_VSS_Mn7@851_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@850 N_OUT7_Mn7@850_d N_OUT6_Mn7@850_g N_VSS_Mn7@850_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@851 N_OUT7_Mp7@851_d N_OUT6_Mp7@851_g N_VDD_Mp7@851_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@850 N_OUT7_Mp7@850_d N_OUT6_Mp7@850_g N_VDD_Mp7@850_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@849 N_OUT7_Mn7@849_d N_OUT6_Mn7@849_g N_VSS_Mn7@849_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@848 N_OUT7_Mn7@848_d N_OUT6_Mn7@848_g N_VSS_Mn7@848_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@849 N_OUT7_Mp7@849_d N_OUT6_Mp7@849_g N_VDD_Mp7@849_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@848 N_OUT7_Mp7@848_d N_OUT6_Mp7@848_g N_VDD_Mp7@848_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@847 N_OUT7_Mn7@847_d N_OUT6_Mn7@847_g N_VSS_Mn7@847_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@846 N_OUT7_Mn7@846_d N_OUT6_Mn7@846_g N_VSS_Mn7@846_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@847 N_OUT7_Mp7@847_d N_OUT6_Mp7@847_g N_VDD_Mp7@847_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@846 N_OUT7_Mp7@846_d N_OUT6_Mp7@846_g N_VDD_Mp7@846_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@845 N_OUT7_Mn7@845_d N_OUT6_Mn7@845_g N_VSS_Mn7@845_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@844 N_OUT7_Mn7@844_d N_OUT6_Mn7@844_g N_VSS_Mn7@844_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@845 N_OUT7_Mp7@845_d N_OUT6_Mp7@845_g N_VDD_Mp7@845_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@844 N_OUT7_Mp7@844_d N_OUT6_Mp7@844_g N_VDD_Mp7@844_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@843 N_OUT7_Mn7@843_d N_OUT6_Mn7@843_g N_VSS_Mn7@843_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@842 N_OUT7_Mn7@842_d N_OUT6_Mn7@842_g N_VSS_Mn7@842_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@843 N_OUT7_Mp7@843_d N_OUT6_Mp7@843_g N_VDD_Mp7@843_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@842 N_OUT7_Mp7@842_d N_OUT6_Mp7@842_g N_VDD_Mp7@842_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@841 N_OUT7_Mn7@841_d N_OUT6_Mn7@841_g N_VSS_Mn7@841_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@840 N_OUT7_Mn7@840_d N_OUT6_Mn7@840_g N_VSS_Mn7@840_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@841 N_OUT7_Mp7@841_d N_OUT6_Mp7@841_g N_VDD_Mp7@841_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@840 N_OUT7_Mp7@840_d N_OUT6_Mp7@840_g N_VDD_Mp7@840_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@839 N_OUT7_Mn7@839_d N_OUT6_Mn7@839_g N_VSS_Mn7@839_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@838 N_OUT7_Mn7@838_d N_OUT6_Mn7@838_g N_VSS_Mn7@838_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@839 N_OUT7_Mp7@839_d N_OUT6_Mp7@839_g N_VDD_Mp7@839_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@838 N_OUT7_Mp7@838_d N_OUT6_Mp7@838_g N_VDD_Mp7@838_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@837 N_OUT7_Mn7@837_d N_OUT6_Mn7@837_g N_VSS_Mn7@837_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@836 N_OUT7_Mn7@836_d N_OUT6_Mn7@836_g N_VSS_Mn7@836_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@837 N_OUT7_Mp7@837_d N_OUT6_Mp7@837_g N_VDD_Mp7@837_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@836 N_OUT7_Mp7@836_d N_OUT6_Mp7@836_g N_VDD_Mp7@836_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@835 N_OUT7_Mn7@835_d N_OUT6_Mn7@835_g N_VSS_Mn7@835_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@834 N_OUT7_Mn7@834_d N_OUT6_Mn7@834_g N_VSS_Mn7@834_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@835 N_OUT7_Mp7@835_d N_OUT6_Mp7@835_g N_VDD_Mp7@835_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@834 N_OUT7_Mp7@834_d N_OUT6_Mp7@834_g N_VDD_Mp7@834_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@833 N_OUT7_Mn7@833_d N_OUT6_Mn7@833_g N_VSS_Mn7@833_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@832 N_OUT7_Mn7@832_d N_OUT6_Mn7@832_g N_VSS_Mn7@832_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@833 N_OUT7_Mp7@833_d N_OUT6_Mp7@833_g N_VDD_Mp7@833_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@832 N_OUT7_Mp7@832_d N_OUT6_Mp7@832_g N_VDD_Mp7@832_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@831 N_OUT7_Mn7@831_d N_OUT6_Mn7@831_g N_VSS_Mn7@831_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@830 N_OUT7_Mn7@830_d N_OUT6_Mn7@830_g N_VSS_Mn7@830_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@831 N_OUT7_Mp7@831_d N_OUT6_Mp7@831_g N_VDD_Mp7@831_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@830 N_OUT7_Mp7@830_d N_OUT6_Mp7@830_g N_VDD_Mp7@830_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@829 N_OUT7_Mn7@829_d N_OUT6_Mn7@829_g N_VSS_Mn7@829_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@828 N_OUT7_Mn7@828_d N_OUT6_Mn7@828_g N_VSS_Mn7@828_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@829 N_OUT7_Mp7@829_d N_OUT6_Mp7@829_g N_VDD_Mp7@829_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@828 N_OUT7_Mp7@828_d N_OUT6_Mp7@828_g N_VDD_Mp7@828_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@827 N_OUT7_Mn7@827_d N_OUT6_Mn7@827_g N_VSS_Mn7@827_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@826 N_OUT7_Mn7@826_d N_OUT6_Mn7@826_g N_VSS_Mn7@826_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@827 N_OUT7_Mp7@827_d N_OUT6_Mp7@827_g N_VDD_Mp7@827_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@826 N_OUT7_Mp7@826_d N_OUT6_Mp7@826_g N_VDD_Mp7@826_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@825 N_OUT7_Mn7@825_d N_OUT6_Mn7@825_g N_VSS_Mn7@825_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@824 N_OUT7_Mn7@824_d N_OUT6_Mn7@824_g N_VSS_Mn7@824_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@825 N_OUT7_Mp7@825_d N_OUT6_Mp7@825_g N_VDD_Mp7@825_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@824 N_OUT7_Mp7@824_d N_OUT6_Mp7@824_g N_VDD_Mp7@824_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@823 N_OUT7_Mn7@823_d N_OUT6_Mn7@823_g N_VSS_Mn7@823_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@822 N_OUT7_Mn7@822_d N_OUT6_Mn7@822_g N_VSS_Mn7@822_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@823 N_OUT7_Mp7@823_d N_OUT6_Mp7@823_g N_VDD_Mp7@823_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@822 N_OUT7_Mp7@822_d N_OUT6_Mp7@822_g N_VDD_Mp7@822_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@821 N_OUT7_Mn7@821_d N_OUT6_Mn7@821_g N_VSS_Mn7@821_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@820 N_OUT7_Mn7@820_d N_OUT6_Mn7@820_g N_VSS_Mn7@820_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@821 N_OUT7_Mp7@821_d N_OUT6_Mp7@821_g N_VDD_Mp7@821_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@820 N_OUT7_Mp7@820_d N_OUT6_Mp7@820_g N_VDD_Mp7@820_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@819 N_OUT7_Mn7@819_d N_OUT6_Mn7@819_g N_VSS_Mn7@819_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@818 N_OUT7_Mn7@818_d N_OUT6_Mn7@818_g N_VSS_Mn7@818_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@819 N_OUT7_Mp7@819_d N_OUT6_Mp7@819_g N_VDD_Mp7@819_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@818 N_OUT7_Mp7@818_d N_OUT6_Mp7@818_g N_VDD_Mp7@818_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@817 N_OUT7_Mn7@817_d N_OUT6_Mn7@817_g N_VSS_Mn7@817_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@816 N_OUT7_Mn7@816_d N_OUT6_Mn7@816_g N_VSS_Mn7@816_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@817 N_OUT7_Mp7@817_d N_OUT6_Mp7@817_g N_VDD_Mp7@817_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@816 N_OUT7_Mp7@816_d N_OUT6_Mp7@816_g N_VDD_Mp7@816_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@815 N_OUT7_Mn7@815_d N_OUT6_Mn7@815_g N_VSS_Mn7@815_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@814 N_OUT7_Mn7@814_d N_OUT6_Mn7@814_g N_VSS_Mn7@814_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@815 N_OUT7_Mp7@815_d N_OUT6_Mp7@815_g N_VDD_Mp7@815_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@814 N_OUT7_Mp7@814_d N_OUT6_Mp7@814_g N_VDD_Mp7@814_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@813 N_OUT7_Mn7@813_d N_OUT6_Mn7@813_g N_VSS_Mn7@813_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@812 N_OUT7_Mn7@812_d N_OUT6_Mn7@812_g N_VSS_Mn7@812_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@813 N_OUT7_Mp7@813_d N_OUT6_Mp7@813_g N_VDD_Mp7@813_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@812 N_OUT7_Mp7@812_d N_OUT6_Mp7@812_g N_VDD_Mp7@812_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@811 N_OUT7_Mn7@811_d N_OUT6_Mn7@811_g N_VSS_Mn7@811_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@810 N_OUT7_Mn7@810_d N_OUT6_Mn7@810_g N_VSS_Mn7@810_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@811 N_OUT7_Mp7@811_d N_OUT6_Mp7@811_g N_VDD_Mp7@811_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@810 N_OUT7_Mp7@810_d N_OUT6_Mp7@810_g N_VDD_Mp7@810_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@809 N_OUT7_Mn7@809_d N_OUT6_Mn7@809_g N_VSS_Mn7@809_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@808 N_OUT7_Mn7@808_d N_OUT6_Mn7@808_g N_VSS_Mn7@808_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@809 N_OUT7_Mp7@809_d N_OUT6_Mp7@809_g N_VDD_Mp7@809_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@808 N_OUT7_Mp7@808_d N_OUT6_Mp7@808_g N_VDD_Mp7@808_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@807 N_OUT7_Mn7@807_d N_OUT6_Mn7@807_g N_VSS_Mn7@807_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@806 N_OUT7_Mn7@806_d N_OUT6_Mn7@806_g N_VSS_Mn7@806_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@807 N_OUT7_Mp7@807_d N_OUT6_Mp7@807_g N_VDD_Mp7@807_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@806 N_OUT7_Mp7@806_d N_OUT6_Mp7@806_g N_VDD_Mp7@806_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@805 N_OUT7_Mn7@805_d N_OUT6_Mn7@805_g N_VSS_Mn7@805_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@804 N_OUT7_Mn7@804_d N_OUT6_Mn7@804_g N_VSS_Mn7@804_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@805 N_OUT7_Mp7@805_d N_OUT6_Mp7@805_g N_VDD_Mp7@805_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@804 N_OUT7_Mp7@804_d N_OUT6_Mp7@804_g N_VDD_Mp7@804_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@803 N_OUT7_Mn7@803_d N_OUT6_Mn7@803_g N_VSS_Mn7@803_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@802 N_OUT7_Mn7@802_d N_OUT6_Mn7@802_g N_VSS_Mn7@802_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@803 N_OUT7_Mp7@803_d N_OUT6_Mp7@803_g N_VDD_Mp7@803_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@802 N_OUT7_Mp7@802_d N_OUT6_Mp7@802_g N_VDD_Mp7@802_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@801 N_OUT7_Mn7@801_d N_OUT6_Mn7@801_g N_VSS_Mn7@801_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@800 N_OUT7_Mn7@800_d N_OUT6_Mn7@800_g N_VSS_Mn7@800_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@801 N_OUT7_Mp7@801_d N_OUT6_Mp7@801_g N_VDD_Mp7@801_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@800 N_OUT7_Mp7@800_d N_OUT6_Mp7@800_g N_VDD_Mp7@800_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@799 N_OUT7_Mn7@799_d N_OUT6_Mn7@799_g N_VSS_Mn7@799_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@798 N_OUT7_Mn7@798_d N_OUT6_Mn7@798_g N_VSS_Mn7@798_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@799 N_OUT7_Mp7@799_d N_OUT6_Mp7@799_g N_VDD_Mp7@799_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@798 N_OUT7_Mp7@798_d N_OUT6_Mp7@798_g N_VDD_Mp7@798_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@797 N_OUT7_Mn7@797_d N_OUT6_Mn7@797_g N_VSS_Mn7@797_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@796 N_OUT7_Mn7@796_d N_OUT6_Mn7@796_g N_VSS_Mn7@796_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@797 N_OUT7_Mp7@797_d N_OUT6_Mp7@797_g N_VDD_Mp7@797_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@796 N_OUT7_Mp7@796_d N_OUT6_Mp7@796_g N_VDD_Mp7@796_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@795 N_OUT7_Mn7@795_d N_OUT6_Mn7@795_g N_VSS_Mn7@795_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@794 N_OUT7_Mn7@794_d N_OUT6_Mn7@794_g N_VSS_Mn7@794_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@795 N_OUT7_Mp7@795_d N_OUT6_Mp7@795_g N_VDD_Mp7@795_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@794 N_OUT7_Mp7@794_d N_OUT6_Mp7@794_g N_VDD_Mp7@794_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@793 N_OUT7_Mn7@793_d N_OUT6_Mn7@793_g N_VSS_Mn7@793_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@792 N_OUT7_Mn7@792_d N_OUT6_Mn7@792_g N_VSS_Mn7@792_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@793 N_OUT7_Mp7@793_d N_OUT6_Mp7@793_g N_VDD_Mp7@793_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@792 N_OUT7_Mp7@792_d N_OUT6_Mp7@792_g N_VDD_Mp7@792_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@791 N_OUT7_Mn7@791_d N_OUT6_Mn7@791_g N_VSS_Mn7@791_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@790 N_OUT7_Mn7@790_d N_OUT6_Mn7@790_g N_VSS_Mn7@790_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@791 N_OUT7_Mp7@791_d N_OUT6_Mp7@791_g N_VDD_Mp7@791_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@790 N_OUT7_Mp7@790_d N_OUT6_Mp7@790_g N_VDD_Mp7@790_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@789 N_OUT7_Mn7@789_d N_OUT6_Mn7@789_g N_VSS_Mn7@789_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@788 N_OUT7_Mn7@788_d N_OUT6_Mn7@788_g N_VSS_Mn7@788_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@789 N_OUT7_Mp7@789_d N_OUT6_Mp7@789_g N_VDD_Mp7@789_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@788 N_OUT7_Mp7@788_d N_OUT6_Mp7@788_g N_VDD_Mp7@788_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@787 N_OUT7_Mn7@787_d N_OUT6_Mn7@787_g N_VSS_Mn7@787_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@786 N_OUT7_Mn7@786_d N_OUT6_Mn7@786_g N_VSS_Mn7@786_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@787 N_OUT7_Mp7@787_d N_OUT6_Mp7@787_g N_VDD_Mp7@787_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@786 N_OUT7_Mp7@786_d N_OUT6_Mp7@786_g N_VDD_Mp7@786_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@785 N_OUT7_Mn7@785_d N_OUT6_Mn7@785_g N_VSS_Mn7@785_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@784 N_OUT7_Mn7@784_d N_OUT6_Mn7@784_g N_VSS_Mn7@784_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@785 N_OUT7_Mp7@785_d N_OUT6_Mp7@785_g N_VDD_Mp7@785_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@784 N_OUT7_Mp7@784_d N_OUT6_Mp7@784_g N_VDD_Mp7@784_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@783 N_OUT7_Mn7@783_d N_OUT6_Mn7@783_g N_VSS_Mn7@783_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@782 N_OUT7_Mn7@782_d N_OUT6_Mn7@782_g N_VSS_Mn7@782_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@783 N_OUT7_Mp7@783_d N_OUT6_Mp7@783_g N_VDD_Mp7@783_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@782 N_OUT7_Mp7@782_d N_OUT6_Mp7@782_g N_VDD_Mp7@782_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@781 N_OUT7_Mn7@781_d N_OUT6_Mn7@781_g N_VSS_Mn7@781_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@780 N_OUT7_Mn7@780_d N_OUT6_Mn7@780_g N_VSS_Mn7@780_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@781 N_OUT7_Mp7@781_d N_OUT6_Mp7@781_g N_VDD_Mp7@781_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@780 N_OUT7_Mp7@780_d N_OUT6_Mp7@780_g N_VDD_Mp7@780_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@779 N_OUT7_Mn7@779_d N_OUT6_Mn7@779_g N_VSS_Mn7@779_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@778 N_OUT7_Mn7@778_d N_OUT6_Mn7@778_g N_VSS_Mn7@778_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@779 N_OUT7_Mp7@779_d N_OUT6_Mp7@779_g N_VDD_Mp7@779_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@778 N_OUT7_Mp7@778_d N_OUT6_Mp7@778_g N_VDD_Mp7@778_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@777 N_OUT7_Mn7@777_d N_OUT6_Mn7@777_g N_VSS_Mn7@777_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@776 N_OUT7_Mn7@776_d N_OUT6_Mn7@776_g N_VSS_Mn7@776_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@777 N_OUT7_Mp7@777_d N_OUT6_Mp7@777_g N_VDD_Mp7@777_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@776 N_OUT7_Mp7@776_d N_OUT6_Mp7@776_g N_VDD_Mp7@776_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@775 N_OUT7_Mn7@775_d N_OUT6_Mn7@775_g N_VSS_Mn7@775_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@774 N_OUT7_Mn7@774_d N_OUT6_Mn7@774_g N_VSS_Mn7@774_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@775 N_OUT7_Mp7@775_d N_OUT6_Mp7@775_g N_VDD_Mp7@775_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@774 N_OUT7_Mp7@774_d N_OUT6_Mp7@774_g N_VDD_Mp7@774_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@773 N_OUT7_Mn7@773_d N_OUT6_Mn7@773_g N_VSS_Mn7@773_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@772 N_OUT7_Mn7@772_d N_OUT6_Mn7@772_g N_VSS_Mn7@772_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@773 N_OUT7_Mp7@773_d N_OUT6_Mp7@773_g N_VDD_Mp7@773_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@772 N_OUT7_Mp7@772_d N_OUT6_Mp7@772_g N_VDD_Mp7@772_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@771 N_OUT7_Mn7@771_d N_OUT6_Mn7@771_g N_VSS_Mn7@771_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@770 N_OUT7_Mn7@770_d N_OUT6_Mn7@770_g N_VSS_Mn7@770_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@771 N_OUT7_Mp7@771_d N_OUT6_Mp7@771_g N_VDD_Mp7@771_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@770 N_OUT7_Mp7@770_d N_OUT6_Mp7@770_g N_VDD_Mp7@770_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@769 N_OUT7_Mn7@769_d N_OUT6_Mn7@769_g N_VSS_Mn7@769_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@768 N_OUT7_Mn7@768_d N_OUT6_Mn7@768_g N_VSS_Mn7@768_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@769 N_OUT7_Mp7@769_d N_OUT6_Mp7@769_g N_VDD_Mp7@769_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@768 N_OUT7_Mp7@768_d N_OUT6_Mp7@768_g N_VDD_Mp7@768_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@767 N_OUT7_Mn7@767_d N_OUT6_Mn7@767_g N_VSS_Mn7@767_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@766 N_OUT7_Mn7@766_d N_OUT6_Mn7@766_g N_VSS_Mn7@766_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@767 N_OUT7_Mp7@767_d N_OUT6_Mp7@767_g N_VDD_Mp7@767_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@766 N_OUT7_Mp7@766_d N_OUT6_Mp7@766_g N_VDD_Mp7@766_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@765 N_OUT7_Mn7@765_d N_OUT6_Mn7@765_g N_VSS_Mn7@765_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@764 N_OUT7_Mn7@764_d N_OUT6_Mn7@764_g N_VSS_Mn7@764_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@765 N_OUT7_Mp7@765_d N_OUT6_Mp7@765_g N_VDD_Mp7@765_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@764 N_OUT7_Mp7@764_d N_OUT6_Mp7@764_g N_VDD_Mp7@764_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@763 N_OUT7_Mn7@763_d N_OUT6_Mn7@763_g N_VSS_Mn7@763_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@762 N_OUT7_Mn7@762_d N_OUT6_Mn7@762_g N_VSS_Mn7@762_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@763 N_OUT7_Mp7@763_d N_OUT6_Mp7@763_g N_VDD_Mp7@763_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@762 N_OUT7_Mp7@762_d N_OUT6_Mp7@762_g N_VDD_Mp7@762_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@761 N_OUT7_Mn7@761_d N_OUT6_Mn7@761_g N_VSS_Mn7@761_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@760 N_OUT7_Mn7@760_d N_OUT6_Mn7@760_g N_VSS_Mn7@760_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@761 N_OUT7_Mp7@761_d N_OUT6_Mp7@761_g N_VDD_Mp7@761_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@760 N_OUT7_Mp7@760_d N_OUT6_Mp7@760_g N_VDD_Mp7@760_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@759 N_OUT7_Mn7@759_d N_OUT6_Mn7@759_g N_VSS_Mn7@759_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@758 N_OUT7_Mn7@758_d N_OUT6_Mn7@758_g N_VSS_Mn7@758_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@759 N_OUT7_Mp7@759_d N_OUT6_Mp7@759_g N_VDD_Mp7@759_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@758 N_OUT7_Mp7@758_d N_OUT6_Mp7@758_g N_VDD_Mp7@758_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@757 N_OUT7_Mn7@757_d N_OUT6_Mn7@757_g N_VSS_Mn7@757_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@756 N_OUT7_Mn7@756_d N_OUT6_Mn7@756_g N_VSS_Mn7@756_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@757 N_OUT7_Mp7@757_d N_OUT6_Mp7@757_g N_VDD_Mp7@757_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@756 N_OUT7_Mp7@756_d N_OUT6_Mp7@756_g N_VDD_Mp7@756_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@755 N_OUT7_Mn7@755_d N_OUT6_Mn7@755_g N_VSS_Mn7@755_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@754 N_OUT7_Mn7@754_d N_OUT6_Mn7@754_g N_VSS_Mn7@754_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@755 N_OUT7_Mp7@755_d N_OUT6_Mp7@755_g N_VDD_Mp7@755_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@754 N_OUT7_Mp7@754_d N_OUT6_Mp7@754_g N_VDD_Mp7@754_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@753 N_OUT7_Mn7@753_d N_OUT6_Mn7@753_g N_VSS_Mn7@753_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@752 N_OUT7_Mn7@752_d N_OUT6_Mn7@752_g N_VSS_Mn7@752_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@753 N_OUT7_Mp7@753_d N_OUT6_Mp7@753_g N_VDD_Mp7@753_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@752 N_OUT7_Mp7@752_d N_OUT6_Mp7@752_g N_VDD_Mp7@752_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@751 N_OUT7_Mn7@751_d N_OUT6_Mn7@751_g N_VSS_Mn7@751_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@750 N_OUT7_Mn7@750_d N_OUT6_Mn7@750_g N_VSS_Mn7@750_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@751 N_OUT7_Mp7@751_d N_OUT6_Mp7@751_g N_VDD_Mp7@751_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@750 N_OUT7_Mp7@750_d N_OUT6_Mp7@750_g N_VDD_Mp7@750_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@749 N_OUT7_Mn7@749_d N_OUT6_Mn7@749_g N_VSS_Mn7@749_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@748 N_OUT7_Mn7@748_d N_OUT6_Mn7@748_g N_VSS_Mn7@748_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@749 N_OUT7_Mp7@749_d N_OUT6_Mp7@749_g N_VDD_Mp7@749_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@748 N_OUT7_Mp7@748_d N_OUT6_Mp7@748_g N_VDD_Mp7@748_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@747 N_OUT7_Mn7@747_d N_OUT6_Mn7@747_g N_VSS_Mn7@747_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@746 N_OUT7_Mn7@746_d N_OUT6_Mn7@746_g N_VSS_Mn7@746_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@747 N_OUT7_Mp7@747_d N_OUT6_Mp7@747_g N_VDD_Mp7@747_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@746 N_OUT7_Mp7@746_d N_OUT6_Mp7@746_g N_VDD_Mp7@746_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@745 N_OUT7_Mn7@745_d N_OUT6_Mn7@745_g N_VSS_Mn7@745_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@744 N_OUT7_Mn7@744_d N_OUT6_Mn7@744_g N_VSS_Mn7@744_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@745 N_OUT7_Mp7@745_d N_OUT6_Mp7@745_g N_VDD_Mp7@745_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@744 N_OUT7_Mp7@744_d N_OUT6_Mp7@744_g N_VDD_Mp7@744_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@743 N_OUT7_Mn7@743_d N_OUT6_Mn7@743_g N_VSS_Mn7@743_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@742 N_OUT7_Mn7@742_d N_OUT6_Mn7@742_g N_VSS_Mn7@742_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@743 N_OUT7_Mp7@743_d N_OUT6_Mp7@743_g N_VDD_Mp7@743_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@742 N_OUT7_Mp7@742_d N_OUT6_Mp7@742_g N_VDD_Mp7@742_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@741 N_OUT7_Mn7@741_d N_OUT6_Mn7@741_g N_VSS_Mn7@741_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@740 N_OUT7_Mn7@740_d N_OUT6_Mn7@740_g N_VSS_Mn7@740_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@741 N_OUT7_Mp7@741_d N_OUT6_Mp7@741_g N_VDD_Mp7@741_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@740 N_OUT7_Mp7@740_d N_OUT6_Mp7@740_g N_VDD_Mp7@740_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@739 N_OUT7_Mn7@739_d N_OUT6_Mn7@739_g N_VSS_Mn7@739_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@738 N_OUT7_Mn7@738_d N_OUT6_Mn7@738_g N_VSS_Mn7@738_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@739 N_OUT7_Mp7@739_d N_OUT6_Mp7@739_g N_VDD_Mp7@739_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@738 N_OUT7_Mp7@738_d N_OUT6_Mp7@738_g N_VDD_Mp7@738_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@737 N_OUT7_Mn7@737_d N_OUT6_Mn7@737_g N_VSS_Mn7@737_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@736 N_OUT7_Mn7@736_d N_OUT6_Mn7@736_g N_VSS_Mn7@736_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@737 N_OUT7_Mp7@737_d N_OUT6_Mp7@737_g N_VDD_Mp7@737_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@736 N_OUT7_Mp7@736_d N_OUT6_Mp7@736_g N_VDD_Mp7@736_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@735 N_OUT7_Mn7@735_d N_OUT6_Mn7@735_g N_VSS_Mn7@735_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@734 N_OUT7_Mn7@734_d N_OUT6_Mn7@734_g N_VSS_Mn7@734_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@735 N_OUT7_Mp7@735_d N_OUT6_Mp7@735_g N_VDD_Mp7@735_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@734 N_OUT7_Mp7@734_d N_OUT6_Mp7@734_g N_VDD_Mp7@734_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@733 N_OUT7_Mn7@733_d N_OUT6_Mn7@733_g N_VSS_Mn7@733_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@732 N_OUT7_Mn7@732_d N_OUT6_Mn7@732_g N_VSS_Mn7@732_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@733 N_OUT7_Mp7@733_d N_OUT6_Mp7@733_g N_VDD_Mp7@733_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@732 N_OUT7_Mp7@732_d N_OUT6_Mp7@732_g N_VDD_Mp7@732_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@731 N_OUT7_Mn7@731_d N_OUT6_Mn7@731_g N_VSS_Mn7@731_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@730 N_OUT7_Mn7@730_d N_OUT6_Mn7@730_g N_VSS_Mn7@730_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@731 N_OUT7_Mp7@731_d N_OUT6_Mp7@731_g N_VDD_Mp7@731_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@730 N_OUT7_Mp7@730_d N_OUT6_Mp7@730_g N_VDD_Mp7@730_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@729 N_OUT7_Mn7@729_d N_OUT6_Mn7@729_g N_VSS_Mn7@729_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@728 N_OUT7_Mn7@728_d N_OUT6_Mn7@728_g N_VSS_Mn7@728_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@729 N_OUT7_Mp7@729_d N_OUT6_Mp7@729_g N_VDD_Mp7@729_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@728 N_OUT7_Mp7@728_d N_OUT6_Mp7@728_g N_VDD_Mp7@728_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@727 N_OUT7_Mn7@727_d N_OUT6_Mn7@727_g N_VSS_Mn7@727_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@726 N_OUT7_Mn7@726_d N_OUT6_Mn7@726_g N_VSS_Mn7@726_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@727 N_OUT7_Mp7@727_d N_OUT6_Mp7@727_g N_VDD_Mp7@727_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@726 N_OUT7_Mp7@726_d N_OUT6_Mp7@726_g N_VDD_Mp7@726_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@725 N_OUT7_Mn7@725_d N_OUT6_Mn7@725_g N_VSS_Mn7@725_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@724 N_OUT7_Mn7@724_d N_OUT6_Mn7@724_g N_VSS_Mn7@724_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@725 N_OUT7_Mp7@725_d N_OUT6_Mp7@725_g N_VDD_Mp7@725_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@724 N_OUT7_Mp7@724_d N_OUT6_Mp7@724_g N_VDD_Mp7@724_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@723 N_OUT7_Mn7@723_d N_OUT6_Mn7@723_g N_VSS_Mn7@723_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@722 N_OUT7_Mn7@722_d N_OUT6_Mn7@722_g N_VSS_Mn7@722_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@723 N_OUT7_Mp7@723_d N_OUT6_Mp7@723_g N_VDD_Mp7@723_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@722 N_OUT7_Mp7@722_d N_OUT6_Mp7@722_g N_VDD_Mp7@722_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@721 N_OUT7_Mn7@721_d N_OUT6_Mn7@721_g N_VSS_Mn7@721_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@720 N_OUT7_Mn7@720_d N_OUT6_Mn7@720_g N_VSS_Mn7@720_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@721 N_OUT7_Mp7@721_d N_OUT6_Mp7@721_g N_VDD_Mp7@721_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@720 N_OUT7_Mp7@720_d N_OUT6_Mp7@720_g N_VDD_Mp7@720_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@719 N_OUT7_Mn7@719_d N_OUT6_Mn7@719_g N_VSS_Mn7@719_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@718 N_OUT7_Mn7@718_d N_OUT6_Mn7@718_g N_VSS_Mn7@718_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@719 N_OUT7_Mp7@719_d N_OUT6_Mp7@719_g N_VDD_Mp7@719_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@718 N_OUT7_Mp7@718_d N_OUT6_Mp7@718_g N_VDD_Mp7@718_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@717 N_OUT7_Mn7@717_d N_OUT6_Mn7@717_g N_VSS_Mn7@717_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@716 N_OUT7_Mn7@716_d N_OUT6_Mn7@716_g N_VSS_Mn7@716_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@717 N_OUT7_Mp7@717_d N_OUT6_Mp7@717_g N_VDD_Mp7@717_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@716 N_OUT7_Mp7@716_d N_OUT6_Mp7@716_g N_VDD_Mp7@716_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@715 N_OUT7_Mn7@715_d N_OUT6_Mn7@715_g N_VSS_Mn7@715_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@714 N_OUT7_Mn7@714_d N_OUT6_Mn7@714_g N_VSS_Mn7@714_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@715 N_OUT7_Mp7@715_d N_OUT6_Mp7@715_g N_VDD_Mp7@715_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@714 N_OUT7_Mp7@714_d N_OUT6_Mp7@714_g N_VDD_Mp7@714_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@713 N_OUT7_Mn7@713_d N_OUT6_Mn7@713_g N_VSS_Mn7@713_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@712 N_OUT7_Mn7@712_d N_OUT6_Mn7@712_g N_VSS_Mn7@712_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@713 N_OUT7_Mp7@713_d N_OUT6_Mp7@713_g N_VDD_Mp7@713_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@712 N_OUT7_Mp7@712_d N_OUT6_Mp7@712_g N_VDD_Mp7@712_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@711 N_OUT7_Mn7@711_d N_OUT6_Mn7@711_g N_VSS_Mn7@711_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@710 N_OUT7_Mn7@710_d N_OUT6_Mn7@710_g N_VSS_Mn7@710_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@711 N_OUT7_Mp7@711_d N_OUT6_Mp7@711_g N_VDD_Mp7@711_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@710 N_OUT7_Mp7@710_d N_OUT6_Mp7@710_g N_VDD_Mp7@710_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@709 N_OUT7_Mn7@709_d N_OUT6_Mn7@709_g N_VSS_Mn7@709_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@708 N_OUT7_Mn7@708_d N_OUT6_Mn7@708_g N_VSS_Mn7@708_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@709 N_OUT7_Mp7@709_d N_OUT6_Mp7@709_g N_VDD_Mp7@709_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@708 N_OUT7_Mp7@708_d N_OUT6_Mp7@708_g N_VDD_Mp7@708_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@707 N_OUT7_Mn7@707_d N_OUT6_Mn7@707_g N_VSS_Mn7@707_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@706 N_OUT7_Mn7@706_d N_OUT6_Mn7@706_g N_VSS_Mn7@706_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@707 N_OUT7_Mp7@707_d N_OUT6_Mp7@707_g N_VDD_Mp7@707_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@706 N_OUT7_Mp7@706_d N_OUT6_Mp7@706_g N_VDD_Mp7@706_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@705 N_OUT7_Mn7@705_d N_OUT6_Mn7@705_g N_VSS_Mn7@705_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@704 N_OUT7_Mn7@704_d N_OUT6_Mn7@704_g N_VSS_Mn7@704_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@705 N_OUT7_Mp7@705_d N_OUT6_Mp7@705_g N_VDD_Mp7@705_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@704 N_OUT7_Mp7@704_d N_OUT6_Mp7@704_g N_VDD_Mp7@704_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@703 N_OUT7_Mn7@703_d N_OUT6_Mn7@703_g N_VSS_Mn7@703_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@702 N_OUT7_Mn7@702_d N_OUT6_Mn7@702_g N_VSS_Mn7@702_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@703 N_OUT7_Mp7@703_d N_OUT6_Mp7@703_g N_VDD_Mp7@703_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@702 N_OUT7_Mp7@702_d N_OUT6_Mp7@702_g N_VDD_Mp7@702_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@701 N_OUT7_Mn7@701_d N_OUT6_Mn7@701_g N_VSS_Mn7@701_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@700 N_OUT7_Mn7@700_d N_OUT6_Mn7@700_g N_VSS_Mn7@700_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@701 N_OUT7_Mp7@701_d N_OUT6_Mp7@701_g N_VDD_Mp7@701_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@700 N_OUT7_Mp7@700_d N_OUT6_Mp7@700_g N_VDD_Mp7@700_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@699 N_OUT7_Mn7@699_d N_OUT6_Mn7@699_g N_VSS_Mn7@699_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@698 N_OUT7_Mn7@698_d N_OUT6_Mn7@698_g N_VSS_Mn7@698_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@699 N_OUT7_Mp7@699_d N_OUT6_Mp7@699_g N_VDD_Mp7@699_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@698 N_OUT7_Mp7@698_d N_OUT6_Mp7@698_g N_VDD_Mp7@698_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@697 N_OUT7_Mn7@697_d N_OUT6_Mn7@697_g N_VSS_Mn7@697_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@696 N_OUT7_Mn7@696_d N_OUT6_Mn7@696_g N_VSS_Mn7@696_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@697 N_OUT7_Mp7@697_d N_OUT6_Mp7@697_g N_VDD_Mp7@697_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@696 N_OUT7_Mp7@696_d N_OUT6_Mp7@696_g N_VDD_Mp7@696_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@695 N_OUT7_Mn7@695_d N_OUT6_Mn7@695_g N_VSS_Mn7@695_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@694 N_OUT7_Mn7@694_d N_OUT6_Mn7@694_g N_VSS_Mn7@694_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@695 N_OUT7_Mp7@695_d N_OUT6_Mp7@695_g N_VDD_Mp7@695_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@694 N_OUT7_Mp7@694_d N_OUT6_Mp7@694_g N_VDD_Mp7@694_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@693 N_OUT7_Mn7@693_d N_OUT6_Mn7@693_g N_VSS_Mn7@693_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@692 N_OUT7_Mn7@692_d N_OUT6_Mn7@692_g N_VSS_Mn7@692_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@693 N_OUT7_Mp7@693_d N_OUT6_Mp7@693_g N_VDD_Mp7@693_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@692 N_OUT7_Mp7@692_d N_OUT6_Mp7@692_g N_VDD_Mp7@692_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@691 N_OUT7_Mn7@691_d N_OUT6_Mn7@691_g N_VSS_Mn7@691_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@690 N_OUT7_Mn7@690_d N_OUT6_Mn7@690_g N_VSS_Mn7@690_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@691 N_OUT7_Mp7@691_d N_OUT6_Mp7@691_g N_VDD_Mp7@691_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@690 N_OUT7_Mp7@690_d N_OUT6_Mp7@690_g N_VDD_Mp7@690_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@689 N_OUT7_Mn7@689_d N_OUT6_Mn7@689_g N_VSS_Mn7@689_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@688 N_OUT7_Mn7@688_d N_OUT6_Mn7@688_g N_VSS_Mn7@688_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@689 N_OUT7_Mp7@689_d N_OUT6_Mp7@689_g N_VDD_Mp7@689_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@688 N_OUT7_Mp7@688_d N_OUT6_Mp7@688_g N_VDD_Mp7@688_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@687 N_OUT7_Mn7@687_d N_OUT6_Mn7@687_g N_VSS_Mn7@687_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@686 N_OUT7_Mn7@686_d N_OUT6_Mn7@686_g N_VSS_Mn7@686_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@687 N_OUT7_Mp7@687_d N_OUT6_Mp7@687_g N_VDD_Mp7@687_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@686 N_OUT7_Mp7@686_d N_OUT6_Mp7@686_g N_VDD_Mp7@686_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@685 N_OUT7_Mn7@685_d N_OUT6_Mn7@685_g N_VSS_Mn7@685_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@684 N_OUT7_Mn7@684_d N_OUT6_Mn7@684_g N_VSS_Mn7@684_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@685 N_OUT7_Mp7@685_d N_OUT6_Mp7@685_g N_VDD_Mp7@685_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@684 N_OUT7_Mp7@684_d N_OUT6_Mp7@684_g N_VDD_Mp7@684_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@683 N_OUT7_Mn7@683_d N_OUT6_Mn7@683_g N_VSS_Mn7@683_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@682 N_OUT7_Mn7@682_d N_OUT6_Mn7@682_g N_VSS_Mn7@682_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@683 N_OUT7_Mp7@683_d N_OUT6_Mp7@683_g N_VDD_Mp7@683_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@682 N_OUT7_Mp7@682_d N_OUT6_Mp7@682_g N_VDD_Mp7@682_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@681 N_OUT7_Mn7@681_d N_OUT6_Mn7@681_g N_VSS_Mn7@681_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@680 N_OUT7_Mn7@680_d N_OUT6_Mn7@680_g N_VSS_Mn7@680_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@681 N_OUT7_Mp7@681_d N_OUT6_Mp7@681_g N_VDD_Mp7@681_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@680 N_OUT7_Mp7@680_d N_OUT6_Mp7@680_g N_VDD_Mp7@680_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@679 N_OUT7_Mn7@679_d N_OUT6_Mn7@679_g N_VSS_Mn7@679_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@678 N_OUT7_Mn7@678_d N_OUT6_Mn7@678_g N_VSS_Mn7@678_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@679 N_OUT7_Mp7@679_d N_OUT6_Mp7@679_g N_VDD_Mp7@679_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@678 N_OUT7_Mp7@678_d N_OUT6_Mp7@678_g N_VDD_Mp7@678_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@677 N_OUT7_Mn7@677_d N_OUT6_Mn7@677_g N_VSS_Mn7@677_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@676 N_OUT7_Mn7@676_d N_OUT6_Mn7@676_g N_VSS_Mn7@676_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@677 N_OUT7_Mp7@677_d N_OUT6_Mp7@677_g N_VDD_Mp7@677_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@676 N_OUT7_Mp7@676_d N_OUT6_Mp7@676_g N_VDD_Mp7@676_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@675 N_OUT7_Mn7@675_d N_OUT6_Mn7@675_g N_VSS_Mn7@675_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@674 N_OUT7_Mn7@674_d N_OUT6_Mn7@674_g N_VSS_Mn7@674_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@675 N_OUT7_Mp7@675_d N_OUT6_Mp7@675_g N_VDD_Mp7@675_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@674 N_OUT7_Mp7@674_d N_OUT6_Mp7@674_g N_VDD_Mp7@674_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@673 N_OUT7_Mn7@673_d N_OUT6_Mn7@673_g N_VSS_Mn7@673_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@672 N_OUT7_Mn7@672_d N_OUT6_Mn7@672_g N_VSS_Mn7@672_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@673 N_OUT7_Mp7@673_d N_OUT6_Mp7@673_g N_VDD_Mp7@673_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@672 N_OUT7_Mp7@672_d N_OUT6_Mp7@672_g N_VDD_Mp7@672_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@671 N_OUT7_Mn7@671_d N_OUT6_Mn7@671_g N_VSS_Mn7@671_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@670 N_OUT7_Mn7@670_d N_OUT6_Mn7@670_g N_VSS_Mn7@670_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@671 N_OUT7_Mp7@671_d N_OUT6_Mp7@671_g N_VDD_Mp7@671_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@670 N_OUT7_Mp7@670_d N_OUT6_Mp7@670_g N_VDD_Mp7@670_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@669 N_OUT7_Mn7@669_d N_OUT6_Mn7@669_g N_VSS_Mn7@669_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@668 N_OUT7_Mn7@668_d N_OUT6_Mn7@668_g N_VSS_Mn7@668_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@669 N_OUT7_Mp7@669_d N_OUT6_Mp7@669_g N_VDD_Mp7@669_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@668 N_OUT7_Mp7@668_d N_OUT6_Mp7@668_g N_VDD_Mp7@668_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@667 N_OUT7_Mn7@667_d N_OUT6_Mn7@667_g N_VSS_Mn7@667_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@666 N_OUT7_Mn7@666_d N_OUT6_Mn7@666_g N_VSS_Mn7@666_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@667 N_OUT7_Mp7@667_d N_OUT6_Mp7@667_g N_VDD_Mp7@667_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@666 N_OUT7_Mp7@666_d N_OUT6_Mp7@666_g N_VDD_Mp7@666_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@665 N_OUT7_Mn7@665_d N_OUT6_Mn7@665_g N_VSS_Mn7@665_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@664 N_OUT7_Mn7@664_d N_OUT6_Mn7@664_g N_VSS_Mn7@664_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@665 N_OUT7_Mp7@665_d N_OUT6_Mp7@665_g N_VDD_Mp7@665_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@664 N_OUT7_Mp7@664_d N_OUT6_Mp7@664_g N_VDD_Mp7@664_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@663 N_OUT7_Mn7@663_d N_OUT6_Mn7@663_g N_VSS_Mn7@663_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@662 N_OUT7_Mn7@662_d N_OUT6_Mn7@662_g N_VSS_Mn7@662_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@663 N_OUT7_Mp7@663_d N_OUT6_Mp7@663_g N_VDD_Mp7@663_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@662 N_OUT7_Mp7@662_d N_OUT6_Mp7@662_g N_VDD_Mp7@662_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@661 N_OUT7_Mn7@661_d N_OUT6_Mn7@661_g N_VSS_Mn7@661_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@660 N_OUT7_Mn7@660_d N_OUT6_Mn7@660_g N_VSS_Mn7@660_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@661 N_OUT7_Mp7@661_d N_OUT6_Mp7@661_g N_VDD_Mp7@661_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@660 N_OUT7_Mp7@660_d N_OUT6_Mp7@660_g N_VDD_Mp7@660_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@659 N_OUT7_Mn7@659_d N_OUT6_Mn7@659_g N_VSS_Mn7@659_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@658 N_OUT7_Mn7@658_d N_OUT6_Mn7@658_g N_VSS_Mn7@658_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@659 N_OUT7_Mp7@659_d N_OUT6_Mp7@659_g N_VDD_Mp7@659_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@658 N_OUT7_Mp7@658_d N_OUT6_Mp7@658_g N_VDD_Mp7@658_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@657 N_OUT7_Mn7@657_d N_OUT6_Mn7@657_g N_VSS_Mn7@657_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@656 N_OUT7_Mn7@656_d N_OUT6_Mn7@656_g N_VSS_Mn7@656_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@657 N_OUT7_Mp7@657_d N_OUT6_Mp7@657_g N_VDD_Mp7@657_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@656 N_OUT7_Mp7@656_d N_OUT6_Mp7@656_g N_VDD_Mp7@656_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@655 N_OUT7_Mn7@655_d N_OUT6_Mn7@655_g N_VSS_Mn7@655_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@654 N_OUT7_Mn7@654_d N_OUT6_Mn7@654_g N_VSS_Mn7@654_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@655 N_OUT7_Mp7@655_d N_OUT6_Mp7@655_g N_VDD_Mp7@655_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@654 N_OUT7_Mp7@654_d N_OUT6_Mp7@654_g N_VDD_Mp7@654_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@653 N_OUT7_Mn7@653_d N_OUT6_Mn7@653_g N_VSS_Mn7@653_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@652 N_OUT7_Mn7@652_d N_OUT6_Mn7@652_g N_VSS_Mn7@652_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@653 N_OUT7_Mp7@653_d N_OUT6_Mp7@653_g N_VDD_Mp7@653_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@652 N_OUT7_Mp7@652_d N_OUT6_Mp7@652_g N_VDD_Mp7@652_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@651 N_OUT7_Mn7@651_d N_OUT6_Mn7@651_g N_VSS_Mn7@651_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@650 N_OUT7_Mn7@650_d N_OUT6_Mn7@650_g N_VSS_Mn7@650_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@651 N_OUT7_Mp7@651_d N_OUT6_Mp7@651_g N_VDD_Mp7@651_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@650 N_OUT7_Mp7@650_d N_OUT6_Mp7@650_g N_VDD_Mp7@650_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@649 N_OUT7_Mn7@649_d N_OUT6_Mn7@649_g N_VSS_Mn7@649_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@648 N_OUT7_Mn7@648_d N_OUT6_Mn7@648_g N_VSS_Mn7@648_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@649 N_OUT7_Mp7@649_d N_OUT6_Mp7@649_g N_VDD_Mp7@649_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@648 N_OUT7_Mp7@648_d N_OUT6_Mp7@648_g N_VDD_Mp7@648_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@647 N_OUT7_Mn7@647_d N_OUT6_Mn7@647_g N_VSS_Mn7@647_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@646 N_OUT7_Mn7@646_d N_OUT6_Mn7@646_g N_VSS_Mn7@646_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@647 N_OUT7_Mp7@647_d N_OUT6_Mp7@647_g N_VDD_Mp7@647_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@646 N_OUT7_Mp7@646_d N_OUT6_Mp7@646_g N_VDD_Mp7@646_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@645 N_OUT7_Mn7@645_d N_OUT6_Mn7@645_g N_VSS_Mn7@645_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@644 N_OUT7_Mn7@644_d N_OUT6_Mn7@644_g N_VSS_Mn7@644_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@645 N_OUT7_Mp7@645_d N_OUT6_Mp7@645_g N_VDD_Mp7@645_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@644 N_OUT7_Mp7@644_d N_OUT6_Mp7@644_g N_VDD_Mp7@644_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@643 N_OUT7_Mn7@643_d N_OUT6_Mn7@643_g N_VSS_Mn7@643_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@642 N_OUT7_Mn7@642_d N_OUT6_Mn7@642_g N_VSS_Mn7@642_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@643 N_OUT7_Mp7@643_d N_OUT6_Mp7@643_g N_VDD_Mp7@643_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@642 N_OUT7_Mp7@642_d N_OUT6_Mp7@642_g N_VDD_Mp7@642_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@641 N_OUT7_Mn7@641_d N_OUT6_Mn7@641_g N_VSS_Mn7@641_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@640 N_OUT7_Mn7@640_d N_OUT6_Mn7@640_g N_VSS_Mn7@640_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@641 N_OUT7_Mp7@641_d N_OUT6_Mp7@641_g N_VDD_Mp7@641_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@640 N_OUT7_Mp7@640_d N_OUT6_Mp7@640_g N_VDD_Mp7@640_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@639 N_OUT7_Mn7@639_d N_OUT6_Mn7@639_g N_VSS_Mn7@639_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@638 N_OUT7_Mn7@638_d N_OUT6_Mn7@638_g N_VSS_Mn7@638_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@639 N_OUT7_Mp7@639_d N_OUT6_Mp7@639_g N_VDD_Mp7@639_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@638 N_OUT7_Mp7@638_d N_OUT6_Mp7@638_g N_VDD_Mp7@638_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@637 N_OUT7_Mn7@637_d N_OUT6_Mn7@637_g N_VSS_Mn7@637_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@636 N_OUT7_Mn7@636_d N_OUT6_Mn7@636_g N_VSS_Mn7@636_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@637 N_OUT7_Mp7@637_d N_OUT6_Mp7@637_g N_VDD_Mp7@637_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@636 N_OUT7_Mp7@636_d N_OUT6_Mp7@636_g N_VDD_Mp7@636_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@635 N_OUT7_Mn7@635_d N_OUT6_Mn7@635_g N_VSS_Mn7@635_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@634 N_OUT7_Mn7@634_d N_OUT6_Mn7@634_g N_VSS_Mn7@634_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@635 N_OUT7_Mp7@635_d N_OUT6_Mp7@635_g N_VDD_Mp7@635_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@634 N_OUT7_Mp7@634_d N_OUT6_Mp7@634_g N_VDD_Mp7@634_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@633 N_OUT7_Mn7@633_d N_OUT6_Mn7@633_g N_VSS_Mn7@633_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@632 N_OUT7_Mn7@632_d N_OUT6_Mn7@632_g N_VSS_Mn7@632_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@633 N_OUT7_Mp7@633_d N_OUT6_Mp7@633_g N_VDD_Mp7@633_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@632 N_OUT7_Mp7@632_d N_OUT6_Mp7@632_g N_VDD_Mp7@632_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@631 N_OUT7_Mn7@631_d N_OUT6_Mn7@631_g N_VSS_Mn7@631_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@630 N_OUT7_Mn7@630_d N_OUT6_Mn7@630_g N_VSS_Mn7@630_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@631 N_OUT7_Mp7@631_d N_OUT6_Mp7@631_g N_VDD_Mp7@631_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@630 N_OUT7_Mp7@630_d N_OUT6_Mp7@630_g N_VDD_Mp7@630_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@629 N_OUT7_Mn7@629_d N_OUT6_Mn7@629_g N_VSS_Mn7@629_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@628 N_OUT7_Mn7@628_d N_OUT6_Mn7@628_g N_VSS_Mn7@628_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@629 N_OUT7_Mp7@629_d N_OUT6_Mp7@629_g N_VDD_Mp7@629_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@628 N_OUT7_Mp7@628_d N_OUT6_Mp7@628_g N_VDD_Mp7@628_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@627 N_OUT7_Mn7@627_d N_OUT6_Mn7@627_g N_VSS_Mn7@627_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@626 N_OUT7_Mn7@626_d N_OUT6_Mn7@626_g N_VSS_Mn7@626_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@627 N_OUT7_Mp7@627_d N_OUT6_Mp7@627_g N_VDD_Mp7@627_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@626 N_OUT7_Mp7@626_d N_OUT6_Mp7@626_g N_VDD_Mp7@626_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@625 N_OUT7_Mn7@625_d N_OUT6_Mn7@625_g N_VSS_Mn7@625_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@624 N_OUT7_Mn7@624_d N_OUT6_Mn7@624_g N_VSS_Mn7@624_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@625 N_OUT7_Mp7@625_d N_OUT6_Mp7@625_g N_VDD_Mp7@625_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@624 N_OUT7_Mp7@624_d N_OUT6_Mp7@624_g N_VDD_Mp7@624_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@623 N_OUT7_Mn7@623_d N_OUT6_Mn7@623_g N_VSS_Mn7@623_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@622 N_OUT7_Mn7@622_d N_OUT6_Mn7@622_g N_VSS_Mn7@622_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@623 N_OUT7_Mp7@623_d N_OUT6_Mp7@623_g N_VDD_Mp7@623_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@622 N_OUT7_Mp7@622_d N_OUT6_Mp7@622_g N_VDD_Mp7@622_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@621 N_OUT7_Mn7@621_d N_OUT6_Mn7@621_g N_VSS_Mn7@621_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@620 N_OUT7_Mn7@620_d N_OUT6_Mn7@620_g N_VSS_Mn7@620_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@621 N_OUT7_Mp7@621_d N_OUT6_Mp7@621_g N_VDD_Mp7@621_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@620 N_OUT7_Mp7@620_d N_OUT6_Mp7@620_g N_VDD_Mp7@620_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@619 N_OUT7_Mn7@619_d N_OUT6_Mn7@619_g N_VSS_Mn7@619_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@618 N_OUT7_Mn7@618_d N_OUT6_Mn7@618_g N_VSS_Mn7@618_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@619 N_OUT7_Mp7@619_d N_OUT6_Mp7@619_g N_VDD_Mp7@619_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@618 N_OUT7_Mp7@618_d N_OUT6_Mp7@618_g N_VDD_Mp7@618_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@617 N_OUT7_Mn7@617_d N_OUT6_Mn7@617_g N_VSS_Mn7@617_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@616 N_OUT7_Mn7@616_d N_OUT6_Mn7@616_g N_VSS_Mn7@616_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@617 N_OUT7_Mp7@617_d N_OUT6_Mp7@617_g N_VDD_Mp7@617_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@616 N_OUT7_Mp7@616_d N_OUT6_Mp7@616_g N_VDD_Mp7@616_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@615 N_OUT7_Mn7@615_d N_OUT6_Mn7@615_g N_VSS_Mn7@615_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@614 N_OUT7_Mn7@614_d N_OUT6_Mn7@614_g N_VSS_Mn7@614_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@615 N_OUT7_Mp7@615_d N_OUT6_Mp7@615_g N_VDD_Mp7@615_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@614 N_OUT7_Mp7@614_d N_OUT6_Mp7@614_g N_VDD_Mp7@614_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@613 N_OUT7_Mn7@613_d N_OUT6_Mn7@613_g N_VSS_Mn7@613_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@612 N_OUT7_Mn7@612_d N_OUT6_Mn7@612_g N_VSS_Mn7@612_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@613 N_OUT7_Mp7@613_d N_OUT6_Mp7@613_g N_VDD_Mp7@613_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@612 N_OUT7_Mp7@612_d N_OUT6_Mp7@612_g N_VDD_Mp7@612_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@611 N_OUT7_Mn7@611_d N_OUT6_Mn7@611_g N_VSS_Mn7@611_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@610 N_OUT7_Mn7@610_d N_OUT6_Mn7@610_g N_VSS_Mn7@610_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@611 N_OUT7_Mp7@611_d N_OUT6_Mp7@611_g N_VDD_Mp7@611_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@610 N_OUT7_Mp7@610_d N_OUT6_Mp7@610_g N_VDD_Mp7@610_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@609 N_OUT7_Mn7@609_d N_OUT6_Mn7@609_g N_VSS_Mn7@609_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@608 N_OUT7_Mn7@608_d N_OUT6_Mn7@608_g N_VSS_Mn7@608_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@609 N_OUT7_Mp7@609_d N_OUT6_Mp7@609_g N_VDD_Mp7@609_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@608 N_OUT7_Mp7@608_d N_OUT6_Mp7@608_g N_VDD_Mp7@608_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@607 N_OUT7_Mn7@607_d N_OUT6_Mn7@607_g N_VSS_Mn7@607_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@606 N_OUT7_Mn7@606_d N_OUT6_Mn7@606_g N_VSS_Mn7@606_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@607 N_OUT7_Mp7@607_d N_OUT6_Mp7@607_g N_VDD_Mp7@607_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@606 N_OUT7_Mp7@606_d N_OUT6_Mp7@606_g N_VDD_Mp7@606_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@605 N_OUT7_Mn7@605_d N_OUT6_Mn7@605_g N_VSS_Mn7@605_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@604 N_OUT7_Mn7@604_d N_OUT6_Mn7@604_g N_VSS_Mn7@604_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@605 N_OUT7_Mp7@605_d N_OUT6_Mp7@605_g N_VDD_Mp7@605_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@604 N_OUT7_Mp7@604_d N_OUT6_Mp7@604_g N_VDD_Mp7@604_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@603 N_OUT7_Mn7@603_d N_OUT6_Mn7@603_g N_VSS_Mn7@603_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@602 N_OUT7_Mn7@602_d N_OUT6_Mn7@602_g N_VSS_Mn7@602_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@603 N_OUT7_Mp7@603_d N_OUT6_Mp7@603_g N_VDD_Mp7@603_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@602 N_OUT7_Mp7@602_d N_OUT6_Mp7@602_g N_VDD_Mp7@602_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@601 N_OUT7_Mn7@601_d N_OUT6_Mn7@601_g N_VSS_Mn7@601_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@600 N_OUT7_Mn7@600_d N_OUT6_Mn7@600_g N_VSS_Mn7@600_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@601 N_OUT7_Mp7@601_d N_OUT6_Mp7@601_g N_VDD_Mp7@601_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@600 N_OUT7_Mp7@600_d N_OUT6_Mp7@600_g N_VDD_Mp7@600_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@599 N_OUT7_Mn7@599_d N_OUT6_Mn7@599_g N_VSS_Mn7@599_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@598 N_OUT7_Mn7@598_d N_OUT6_Mn7@598_g N_VSS_Mn7@598_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@599 N_OUT7_Mp7@599_d N_OUT6_Mp7@599_g N_VDD_Mp7@599_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@598 N_OUT7_Mp7@598_d N_OUT6_Mp7@598_g N_VDD_Mp7@598_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@597 N_OUT7_Mn7@597_d N_OUT6_Mn7@597_g N_VSS_Mn7@597_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@596 N_OUT7_Mn7@596_d N_OUT6_Mn7@596_g N_VSS_Mn7@596_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@597 N_OUT7_Mp7@597_d N_OUT6_Mp7@597_g N_VDD_Mp7@597_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@596 N_OUT7_Mp7@596_d N_OUT6_Mp7@596_g N_VDD_Mp7@596_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@595 N_OUT7_Mn7@595_d N_OUT6_Mn7@595_g N_VSS_Mn7@595_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@594 N_OUT7_Mn7@594_d N_OUT6_Mn7@594_g N_VSS_Mn7@594_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@595 N_OUT7_Mp7@595_d N_OUT6_Mp7@595_g N_VDD_Mp7@595_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@594 N_OUT7_Mp7@594_d N_OUT6_Mp7@594_g N_VDD_Mp7@594_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@593 N_OUT7_Mn7@593_d N_OUT6_Mn7@593_g N_VSS_Mn7@593_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@592 N_OUT7_Mn7@592_d N_OUT6_Mn7@592_g N_VSS_Mn7@592_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@593 N_OUT7_Mp7@593_d N_OUT6_Mp7@593_g N_VDD_Mp7@593_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@592 N_OUT7_Mp7@592_d N_OUT6_Mp7@592_g N_VDD_Mp7@592_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@591 N_OUT7_Mn7@591_d N_OUT6_Mn7@591_g N_VSS_Mn7@591_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@590 N_OUT7_Mn7@590_d N_OUT6_Mn7@590_g N_VSS_Mn7@590_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@591 N_OUT7_Mp7@591_d N_OUT6_Mp7@591_g N_VDD_Mp7@591_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@590 N_OUT7_Mp7@590_d N_OUT6_Mp7@590_g N_VDD_Mp7@590_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@589 N_OUT7_Mn7@589_d N_OUT6_Mn7@589_g N_VSS_Mn7@589_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@588 N_OUT7_Mn7@588_d N_OUT6_Mn7@588_g N_VSS_Mn7@588_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@589 N_OUT7_Mp7@589_d N_OUT6_Mp7@589_g N_VDD_Mp7@589_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@588 N_OUT7_Mp7@588_d N_OUT6_Mp7@588_g N_VDD_Mp7@588_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@587 N_OUT7_Mn7@587_d N_OUT6_Mn7@587_g N_VSS_Mn7@587_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@586 N_OUT7_Mn7@586_d N_OUT6_Mn7@586_g N_VSS_Mn7@586_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@587 N_OUT7_Mp7@587_d N_OUT6_Mp7@587_g N_VDD_Mp7@587_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@586 N_OUT7_Mp7@586_d N_OUT6_Mp7@586_g N_VDD_Mp7@586_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@585 N_OUT7_Mn7@585_d N_OUT6_Mn7@585_g N_VSS_Mn7@585_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@584 N_OUT7_Mn7@584_d N_OUT6_Mn7@584_g N_VSS_Mn7@584_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@585 N_OUT7_Mp7@585_d N_OUT6_Mp7@585_g N_VDD_Mp7@585_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@584 N_OUT7_Mp7@584_d N_OUT6_Mp7@584_g N_VDD_Mp7@584_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@583 N_OUT7_Mn7@583_d N_OUT6_Mn7@583_g N_VSS_Mn7@583_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@582 N_OUT7_Mn7@582_d N_OUT6_Mn7@582_g N_VSS_Mn7@582_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@583 N_OUT7_Mp7@583_d N_OUT6_Mp7@583_g N_VDD_Mp7@583_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@582 N_OUT7_Mp7@582_d N_OUT6_Mp7@582_g N_VDD_Mp7@582_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@581 N_OUT7_Mn7@581_d N_OUT6_Mn7@581_g N_VSS_Mn7@581_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@580 N_OUT7_Mn7@580_d N_OUT6_Mn7@580_g N_VSS_Mn7@580_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@581 N_OUT7_Mp7@581_d N_OUT6_Mp7@581_g N_VDD_Mp7@581_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@580 N_OUT7_Mp7@580_d N_OUT6_Mp7@580_g N_VDD_Mp7@580_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@579 N_OUT7_Mn7@579_d N_OUT6_Mn7@579_g N_VSS_Mn7@579_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@578 N_OUT7_Mn7@578_d N_OUT6_Mn7@578_g N_VSS_Mn7@578_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@579 N_OUT7_Mp7@579_d N_OUT6_Mp7@579_g N_VDD_Mp7@579_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@578 N_OUT7_Mp7@578_d N_OUT6_Mp7@578_g N_VDD_Mp7@578_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@577 N_OUT7_Mn7@577_d N_OUT6_Mn7@577_g N_VSS_Mn7@577_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@576 N_OUT7_Mn7@576_d N_OUT6_Mn7@576_g N_VSS_Mn7@576_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@577 N_OUT7_Mp7@577_d N_OUT6_Mp7@577_g N_VDD_Mp7@577_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@576 N_OUT7_Mp7@576_d N_OUT6_Mp7@576_g N_VDD_Mp7@576_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@575 N_OUT7_Mn7@575_d N_OUT6_Mn7@575_g N_VSS_Mn7@575_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@574 N_OUT7_Mn7@574_d N_OUT6_Mn7@574_g N_VSS_Mn7@574_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@575 N_OUT7_Mp7@575_d N_OUT6_Mp7@575_g N_VDD_Mp7@575_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@574 N_OUT7_Mp7@574_d N_OUT6_Mp7@574_g N_VDD_Mp7@574_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@573 N_OUT7_Mn7@573_d N_OUT6_Mn7@573_g N_VSS_Mn7@573_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@572 N_OUT7_Mn7@572_d N_OUT6_Mn7@572_g N_VSS_Mn7@572_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@573 N_OUT7_Mp7@573_d N_OUT6_Mp7@573_g N_VDD_Mp7@573_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@572 N_OUT7_Mp7@572_d N_OUT6_Mp7@572_g N_VDD_Mp7@572_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@571 N_OUT7_Mn7@571_d N_OUT6_Mn7@571_g N_VSS_Mn7@571_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@570 N_OUT7_Mn7@570_d N_OUT6_Mn7@570_g N_VSS_Mn7@570_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@571 N_OUT7_Mp7@571_d N_OUT6_Mp7@571_g N_VDD_Mp7@571_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@570 N_OUT7_Mp7@570_d N_OUT6_Mp7@570_g N_VDD_Mp7@570_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@569 N_OUT7_Mn7@569_d N_OUT6_Mn7@569_g N_VSS_Mn7@569_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@568 N_OUT7_Mn7@568_d N_OUT6_Mn7@568_g N_VSS_Mn7@568_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@569 N_OUT7_Mp7@569_d N_OUT6_Mp7@569_g N_VDD_Mp7@569_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@568 N_OUT7_Mp7@568_d N_OUT6_Mp7@568_g N_VDD_Mp7@568_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@567 N_OUT7_Mn7@567_d N_OUT6_Mn7@567_g N_VSS_Mn7@567_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@566 N_OUT7_Mn7@566_d N_OUT6_Mn7@566_g N_VSS_Mn7@566_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@567 N_OUT7_Mp7@567_d N_OUT6_Mp7@567_g N_VDD_Mp7@567_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@566 N_OUT7_Mp7@566_d N_OUT6_Mp7@566_g N_VDD_Mp7@566_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@565 N_OUT7_Mn7@565_d N_OUT6_Mn7@565_g N_VSS_Mn7@565_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@564 N_OUT7_Mn7@564_d N_OUT6_Mn7@564_g N_VSS_Mn7@564_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@565 N_OUT7_Mp7@565_d N_OUT6_Mp7@565_g N_VDD_Mp7@565_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@564 N_OUT7_Mp7@564_d N_OUT6_Mp7@564_g N_VDD_Mp7@564_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@563 N_OUT7_Mn7@563_d N_OUT6_Mn7@563_g N_VSS_Mn7@563_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@562 N_OUT7_Mn7@562_d N_OUT6_Mn7@562_g N_VSS_Mn7@562_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@563 N_OUT7_Mp7@563_d N_OUT6_Mp7@563_g N_VDD_Mp7@563_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@562 N_OUT7_Mp7@562_d N_OUT6_Mp7@562_g N_VDD_Mp7@562_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@561 N_OUT7_Mn7@561_d N_OUT6_Mn7@561_g N_VSS_Mn7@561_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@560 N_OUT7_Mn7@560_d N_OUT6_Mn7@560_g N_VSS_Mn7@560_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@561 N_OUT7_Mp7@561_d N_OUT6_Mp7@561_g N_VDD_Mp7@561_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@560 N_OUT7_Mp7@560_d N_OUT6_Mp7@560_g N_VDD_Mp7@560_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@559 N_OUT7_Mn7@559_d N_OUT6_Mn7@559_g N_VSS_Mn7@559_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@558 N_OUT7_Mn7@558_d N_OUT6_Mn7@558_g N_VSS_Mn7@558_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@559 N_OUT7_Mp7@559_d N_OUT6_Mp7@559_g N_VDD_Mp7@559_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@558 N_OUT7_Mp7@558_d N_OUT6_Mp7@558_g N_VDD_Mp7@558_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@557 N_OUT7_Mn7@557_d N_OUT6_Mn7@557_g N_VSS_Mn7@557_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@556 N_OUT7_Mn7@556_d N_OUT6_Mn7@556_g N_VSS_Mn7@556_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@557 N_OUT7_Mp7@557_d N_OUT6_Mp7@557_g N_VDD_Mp7@557_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@556 N_OUT7_Mp7@556_d N_OUT6_Mp7@556_g N_VDD_Mp7@556_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@555 N_OUT7_Mn7@555_d N_OUT6_Mn7@555_g N_VSS_Mn7@555_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@554 N_OUT7_Mn7@554_d N_OUT6_Mn7@554_g N_VSS_Mn7@554_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@555 N_OUT7_Mp7@555_d N_OUT6_Mp7@555_g N_VDD_Mp7@555_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@554 N_OUT7_Mp7@554_d N_OUT6_Mp7@554_g N_VDD_Mp7@554_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@553 N_OUT7_Mn7@553_d N_OUT6_Mn7@553_g N_VSS_Mn7@553_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@552 N_OUT7_Mn7@552_d N_OUT6_Mn7@552_g N_VSS_Mn7@552_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@553 N_OUT7_Mp7@553_d N_OUT6_Mp7@553_g N_VDD_Mp7@553_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@552 N_OUT7_Mp7@552_d N_OUT6_Mp7@552_g N_VDD_Mp7@552_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@551 N_OUT7_Mn7@551_d N_OUT6_Mn7@551_g N_VSS_Mn7@551_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@550 N_OUT7_Mn7@550_d N_OUT6_Mn7@550_g N_VSS_Mn7@550_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@551 N_OUT7_Mp7@551_d N_OUT6_Mp7@551_g N_VDD_Mp7@551_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@550 N_OUT7_Mp7@550_d N_OUT6_Mp7@550_g N_VDD_Mp7@550_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@549 N_OUT7_Mn7@549_d N_OUT6_Mn7@549_g N_VSS_Mn7@549_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@548 N_OUT7_Mn7@548_d N_OUT6_Mn7@548_g N_VSS_Mn7@548_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@549 N_OUT7_Mp7@549_d N_OUT6_Mp7@549_g N_VDD_Mp7@549_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@548 N_OUT7_Mp7@548_d N_OUT6_Mp7@548_g N_VDD_Mp7@548_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@547 N_OUT7_Mn7@547_d N_OUT6_Mn7@547_g N_VSS_Mn7@547_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@546 N_OUT7_Mn7@546_d N_OUT6_Mn7@546_g N_VSS_Mn7@546_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@547 N_OUT7_Mp7@547_d N_OUT6_Mp7@547_g N_VDD_Mp7@547_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@546 N_OUT7_Mp7@546_d N_OUT6_Mp7@546_g N_VDD_Mp7@546_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@545 N_OUT7_Mn7@545_d N_OUT6_Mn7@545_g N_VSS_Mn7@545_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@544 N_OUT7_Mn7@544_d N_OUT6_Mn7@544_g N_VSS_Mn7@544_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@545 N_OUT7_Mp7@545_d N_OUT6_Mp7@545_g N_VDD_Mp7@545_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@544 N_OUT7_Mp7@544_d N_OUT6_Mp7@544_g N_VDD_Mp7@544_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@543 N_OUT7_Mn7@543_d N_OUT6_Mn7@543_g N_VSS_Mn7@543_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@542 N_OUT7_Mn7@542_d N_OUT6_Mn7@542_g N_VSS_Mn7@542_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@543 N_OUT7_Mp7@543_d N_OUT6_Mp7@543_g N_VDD_Mp7@543_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@542 N_OUT7_Mp7@542_d N_OUT6_Mp7@542_g N_VDD_Mp7@542_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@541 N_OUT7_Mn7@541_d N_OUT6_Mn7@541_g N_VSS_Mn7@541_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@540 N_OUT7_Mn7@540_d N_OUT6_Mn7@540_g N_VSS_Mn7@540_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@541 N_OUT7_Mp7@541_d N_OUT6_Mp7@541_g N_VDD_Mp7@541_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@540 N_OUT7_Mp7@540_d N_OUT6_Mp7@540_g N_VDD_Mp7@540_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@539 N_OUT7_Mn7@539_d N_OUT6_Mn7@539_g N_VSS_Mn7@539_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@538 N_OUT7_Mn7@538_d N_OUT6_Mn7@538_g N_VSS_Mn7@538_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@539 N_OUT7_Mp7@539_d N_OUT6_Mp7@539_g N_VDD_Mp7@539_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@538 N_OUT7_Mp7@538_d N_OUT6_Mp7@538_g N_VDD_Mp7@538_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@537 N_OUT7_Mn7@537_d N_OUT6_Mn7@537_g N_VSS_Mn7@537_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@536 N_OUT7_Mn7@536_d N_OUT6_Mn7@536_g N_VSS_Mn7@536_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@537 N_OUT7_Mp7@537_d N_OUT6_Mp7@537_g N_VDD_Mp7@537_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@536 N_OUT7_Mp7@536_d N_OUT6_Mp7@536_g N_VDD_Mp7@536_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@535 N_OUT7_Mn7@535_d N_OUT6_Mn7@535_g N_VSS_Mn7@535_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@534 N_OUT7_Mn7@534_d N_OUT6_Mn7@534_g N_VSS_Mn7@534_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@535 N_OUT7_Mp7@535_d N_OUT6_Mp7@535_g N_VDD_Mp7@535_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@534 N_OUT7_Mp7@534_d N_OUT6_Mp7@534_g N_VDD_Mp7@534_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@533 N_OUT7_Mn7@533_d N_OUT6_Mn7@533_g N_VSS_Mn7@533_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@532 N_OUT7_Mn7@532_d N_OUT6_Mn7@532_g N_VSS_Mn7@532_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@533 N_OUT7_Mp7@533_d N_OUT6_Mp7@533_g N_VDD_Mp7@533_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@532 N_OUT7_Mp7@532_d N_OUT6_Mp7@532_g N_VDD_Mp7@532_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@531 N_OUT7_Mn7@531_d N_OUT6_Mn7@531_g N_VSS_Mn7@531_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@530 N_OUT7_Mn7@530_d N_OUT6_Mn7@530_g N_VSS_Mn7@530_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@531 N_OUT7_Mp7@531_d N_OUT6_Mp7@531_g N_VDD_Mp7@531_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@530 N_OUT7_Mp7@530_d N_OUT6_Mp7@530_g N_VDD_Mp7@530_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@529 N_OUT7_Mn7@529_d N_OUT6_Mn7@529_g N_VSS_Mn7@529_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@528 N_OUT7_Mn7@528_d N_OUT6_Mn7@528_g N_VSS_Mn7@528_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@529 N_OUT7_Mp7@529_d N_OUT6_Mp7@529_g N_VDD_Mp7@529_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@528 N_OUT7_Mp7@528_d N_OUT6_Mp7@528_g N_VDD_Mp7@528_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@527 N_OUT7_Mn7@527_d N_OUT6_Mn7@527_g N_VSS_Mn7@527_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@526 N_OUT7_Mn7@526_d N_OUT6_Mn7@526_g N_VSS_Mn7@526_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@527 N_OUT7_Mp7@527_d N_OUT6_Mp7@527_g N_VDD_Mp7@527_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@526 N_OUT7_Mp7@526_d N_OUT6_Mp7@526_g N_VDD_Mp7@526_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@525 N_OUT7_Mn7@525_d N_OUT6_Mn7@525_g N_VSS_Mn7@525_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@524 N_OUT7_Mn7@524_d N_OUT6_Mn7@524_g N_VSS_Mn7@524_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@525 N_OUT7_Mp7@525_d N_OUT6_Mp7@525_g N_VDD_Mp7@525_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@524 N_OUT7_Mp7@524_d N_OUT6_Mp7@524_g N_VDD_Mp7@524_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@523 N_OUT7_Mn7@523_d N_OUT6_Mn7@523_g N_VSS_Mn7@523_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@522 N_OUT7_Mn7@522_d N_OUT6_Mn7@522_g N_VSS_Mn7@522_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@523 N_OUT7_Mp7@523_d N_OUT6_Mp7@523_g N_VDD_Mp7@523_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@522 N_OUT7_Mp7@522_d N_OUT6_Mp7@522_g N_VDD_Mp7@522_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@521 N_OUT7_Mn7@521_d N_OUT6_Mn7@521_g N_VSS_Mn7@521_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@520 N_OUT7_Mn7@520_d N_OUT6_Mn7@520_g N_VSS_Mn7@520_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@521 N_OUT7_Mp7@521_d N_OUT6_Mp7@521_g N_VDD_Mp7@521_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@520 N_OUT7_Mp7@520_d N_OUT6_Mp7@520_g N_VDD_Mp7@520_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@519 N_OUT7_Mn7@519_d N_OUT6_Mn7@519_g N_VSS_Mn7@519_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@518 N_OUT7_Mn7@518_d N_OUT6_Mn7@518_g N_VSS_Mn7@518_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@519 N_OUT7_Mp7@519_d N_OUT6_Mp7@519_g N_VDD_Mp7@519_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@518 N_OUT7_Mp7@518_d N_OUT6_Mp7@518_g N_VDD_Mp7@518_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@517 N_OUT7_Mn7@517_d N_OUT6_Mn7@517_g N_VSS_Mn7@517_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@516 N_OUT7_Mn7@516_d N_OUT6_Mn7@516_g N_VSS_Mn7@516_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@517 N_OUT7_Mp7@517_d N_OUT6_Mp7@517_g N_VDD_Mp7@517_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@516 N_OUT7_Mp7@516_d N_OUT6_Mp7@516_g N_VDD_Mp7@516_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@515 N_OUT7_Mn7@515_d N_OUT6_Mn7@515_g N_VSS_Mn7@515_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@514 N_OUT7_Mn7@514_d N_OUT6_Mn7@514_g N_VSS_Mn7@514_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@515 N_OUT7_Mp7@515_d N_OUT6_Mp7@515_g N_VDD_Mp7@515_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@514 N_OUT7_Mp7@514_d N_OUT6_Mp7@514_g N_VDD_Mp7@514_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@513 N_OUT7_Mn7@513_d N_OUT6_Mn7@513_g N_VSS_Mn7@513_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@512 N_OUT7_Mn7@512_d N_OUT6_Mn7@512_g N_VSS_Mn7@512_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@513 N_OUT7_Mp7@513_d N_OUT6_Mp7@513_g N_VDD_Mp7@513_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@512 N_OUT7_Mp7@512_d N_OUT6_Mp7@512_g N_VDD_Mp7@512_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@511 N_OUT7_Mn7@511_d N_OUT6_Mn7@511_g N_VSS_Mn7@511_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@510 N_OUT7_Mn7@510_d N_OUT6_Mn7@510_g N_VSS_Mn7@510_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@511 N_OUT7_Mp7@511_d N_OUT6_Mp7@511_g N_VDD_Mp7@511_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@510 N_OUT7_Mp7@510_d N_OUT6_Mp7@510_g N_VDD_Mp7@510_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@509 N_OUT7_Mn7@509_d N_OUT6_Mn7@509_g N_VSS_Mn7@509_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@508 N_OUT7_Mn7@508_d N_OUT6_Mn7@508_g N_VSS_Mn7@508_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@509 N_OUT7_Mp7@509_d N_OUT6_Mp7@509_g N_VDD_Mp7@509_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@508 N_OUT7_Mp7@508_d N_OUT6_Mp7@508_g N_VDD_Mp7@508_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@507 N_OUT7_Mn7@507_d N_OUT6_Mn7@507_g N_VSS_Mn7@507_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@506 N_OUT7_Mn7@506_d N_OUT6_Mn7@506_g N_VSS_Mn7@506_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@507 N_OUT7_Mp7@507_d N_OUT6_Mp7@507_g N_VDD_Mp7@507_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@506 N_OUT7_Mp7@506_d N_OUT6_Mp7@506_g N_VDD_Mp7@506_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@505 N_OUT7_Mn7@505_d N_OUT6_Mn7@505_g N_VSS_Mn7@505_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@504 N_OUT7_Mn7@504_d N_OUT6_Mn7@504_g N_VSS_Mn7@504_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@505 N_OUT7_Mp7@505_d N_OUT6_Mp7@505_g N_VDD_Mp7@505_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@504 N_OUT7_Mp7@504_d N_OUT6_Mp7@504_g N_VDD_Mp7@504_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@503 N_OUT7_Mn7@503_d N_OUT6_Mn7@503_g N_VSS_Mn7@503_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@502 N_OUT7_Mn7@502_d N_OUT6_Mn7@502_g N_VSS_Mn7@502_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@503 N_OUT7_Mp7@503_d N_OUT6_Mp7@503_g N_VDD_Mp7@503_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@502 N_OUT7_Mp7@502_d N_OUT6_Mp7@502_g N_VDD_Mp7@502_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@501 N_OUT7_Mn7@501_d N_OUT6_Mn7@501_g N_VSS_Mn7@501_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@500 N_OUT7_Mn7@500_d N_OUT6_Mn7@500_g N_VSS_Mn7@500_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@501 N_OUT7_Mp7@501_d N_OUT6_Mp7@501_g N_VDD_Mp7@501_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@500 N_OUT7_Mp7@500_d N_OUT6_Mp7@500_g N_VDD_Mp7@500_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@499 N_OUT7_Mn7@499_d N_OUT6_Mn7@499_g N_VSS_Mn7@499_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@498 N_OUT7_Mn7@498_d N_OUT6_Mn7@498_g N_VSS_Mn7@498_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@499 N_OUT7_Mp7@499_d N_OUT6_Mp7@499_g N_VDD_Mp7@499_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@498 N_OUT7_Mp7@498_d N_OUT6_Mp7@498_g N_VDD_Mp7@498_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@497 N_OUT7_Mn7@497_d N_OUT6_Mn7@497_g N_VSS_Mn7@497_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@496 N_OUT7_Mn7@496_d N_OUT6_Mn7@496_g N_VSS_Mn7@496_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@497 N_OUT7_Mp7@497_d N_OUT6_Mp7@497_g N_VDD_Mp7@497_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@496 N_OUT7_Mp7@496_d N_OUT6_Mp7@496_g N_VDD_Mp7@496_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@495 N_OUT7_Mn7@495_d N_OUT6_Mn7@495_g N_VSS_Mn7@495_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@494 N_OUT7_Mn7@494_d N_OUT6_Mn7@494_g N_VSS_Mn7@494_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@495 N_OUT7_Mp7@495_d N_OUT6_Mp7@495_g N_VDD_Mp7@495_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@494 N_OUT7_Mp7@494_d N_OUT6_Mp7@494_g N_VDD_Mp7@494_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@493 N_OUT7_Mn7@493_d N_OUT6_Mn7@493_g N_VSS_Mn7@493_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@492 N_OUT7_Mn7@492_d N_OUT6_Mn7@492_g N_VSS_Mn7@492_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@493 N_OUT7_Mp7@493_d N_OUT6_Mp7@493_g N_VDD_Mp7@493_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@492 N_OUT7_Mp7@492_d N_OUT6_Mp7@492_g N_VDD_Mp7@492_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@491 N_OUT7_Mn7@491_d N_OUT6_Mn7@491_g N_VSS_Mn7@491_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@490 N_OUT7_Mn7@490_d N_OUT6_Mn7@490_g N_VSS_Mn7@490_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@491 N_OUT7_Mp7@491_d N_OUT6_Mp7@491_g N_VDD_Mp7@491_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@490 N_OUT7_Mp7@490_d N_OUT6_Mp7@490_g N_VDD_Mp7@490_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@489 N_OUT7_Mn7@489_d N_OUT6_Mn7@489_g N_VSS_Mn7@489_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@488 N_OUT7_Mn7@488_d N_OUT6_Mn7@488_g N_VSS_Mn7@488_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@489 N_OUT7_Mp7@489_d N_OUT6_Mp7@489_g N_VDD_Mp7@489_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@488 N_OUT7_Mp7@488_d N_OUT6_Mp7@488_g N_VDD_Mp7@488_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@487 N_OUT7_Mn7@487_d N_OUT6_Mn7@487_g N_VSS_Mn7@487_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@486 N_OUT7_Mn7@486_d N_OUT6_Mn7@486_g N_VSS_Mn7@486_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@487 N_OUT7_Mp7@487_d N_OUT6_Mp7@487_g N_VDD_Mp7@487_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@486 N_OUT7_Mp7@486_d N_OUT6_Mp7@486_g N_VDD_Mp7@486_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@485 N_OUT7_Mn7@485_d N_OUT6_Mn7@485_g N_VSS_Mn7@485_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@484 N_OUT7_Mn7@484_d N_OUT6_Mn7@484_g N_VSS_Mn7@484_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@485 N_OUT7_Mp7@485_d N_OUT6_Mp7@485_g N_VDD_Mp7@485_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@484 N_OUT7_Mp7@484_d N_OUT6_Mp7@484_g N_VDD_Mp7@484_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@483 N_OUT7_Mn7@483_d N_OUT6_Mn7@483_g N_VSS_Mn7@483_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@482 N_OUT7_Mn7@482_d N_OUT6_Mn7@482_g N_VSS_Mn7@482_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@483 N_OUT7_Mp7@483_d N_OUT6_Mp7@483_g N_VDD_Mp7@483_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@482 N_OUT7_Mp7@482_d N_OUT6_Mp7@482_g N_VDD_Mp7@482_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@481 N_OUT7_Mn7@481_d N_OUT6_Mn7@481_g N_VSS_Mn7@481_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@480 N_OUT7_Mn7@480_d N_OUT6_Mn7@480_g N_VSS_Mn7@480_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@481 N_OUT7_Mp7@481_d N_OUT6_Mp7@481_g N_VDD_Mp7@481_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@480 N_OUT7_Mp7@480_d N_OUT6_Mp7@480_g N_VDD_Mp7@480_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@479 N_OUT7_Mn7@479_d N_OUT6_Mn7@479_g N_VSS_Mn7@479_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@478 N_OUT7_Mn7@478_d N_OUT6_Mn7@478_g N_VSS_Mn7@478_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@479 N_OUT7_Mp7@479_d N_OUT6_Mp7@479_g N_VDD_Mp7@479_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@478 N_OUT7_Mp7@478_d N_OUT6_Mp7@478_g N_VDD_Mp7@478_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@477 N_OUT7_Mn7@477_d N_OUT6_Mn7@477_g N_VSS_Mn7@477_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@476 N_OUT7_Mn7@476_d N_OUT6_Mn7@476_g N_VSS_Mn7@476_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@477 N_OUT7_Mp7@477_d N_OUT6_Mp7@477_g N_VDD_Mp7@477_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@476 N_OUT7_Mp7@476_d N_OUT6_Mp7@476_g N_VDD_Mp7@476_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@475 N_OUT7_Mn7@475_d N_OUT6_Mn7@475_g N_VSS_Mn7@475_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@474 N_OUT7_Mn7@474_d N_OUT6_Mn7@474_g N_VSS_Mn7@474_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@475 N_OUT7_Mp7@475_d N_OUT6_Mp7@475_g N_VDD_Mp7@475_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@474 N_OUT7_Mp7@474_d N_OUT6_Mp7@474_g N_VDD_Mp7@474_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@473 N_OUT7_Mn7@473_d N_OUT6_Mn7@473_g N_VSS_Mn7@473_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@472 N_OUT7_Mn7@472_d N_OUT6_Mn7@472_g N_VSS_Mn7@472_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@473 N_OUT7_Mp7@473_d N_OUT6_Mp7@473_g N_VDD_Mp7@473_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@472 N_OUT7_Mp7@472_d N_OUT6_Mp7@472_g N_VDD_Mp7@472_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@471 N_OUT7_Mn7@471_d N_OUT6_Mn7@471_g N_VSS_Mn7@471_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@470 N_OUT7_Mn7@470_d N_OUT6_Mn7@470_g N_VSS_Mn7@470_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@471 N_OUT7_Mp7@471_d N_OUT6_Mp7@471_g N_VDD_Mp7@471_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@470 N_OUT7_Mp7@470_d N_OUT6_Mp7@470_g N_VDD_Mp7@470_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@469 N_OUT7_Mn7@469_d N_OUT6_Mn7@469_g N_VSS_Mn7@469_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@468 N_OUT7_Mn7@468_d N_OUT6_Mn7@468_g N_VSS_Mn7@468_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@469 N_OUT7_Mp7@469_d N_OUT6_Mp7@469_g N_VDD_Mp7@469_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@468 N_OUT7_Mp7@468_d N_OUT6_Mp7@468_g N_VDD_Mp7@468_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@467 N_OUT7_Mn7@467_d N_OUT6_Mn7@467_g N_VSS_Mn7@467_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@466 N_OUT7_Mn7@466_d N_OUT6_Mn7@466_g N_VSS_Mn7@466_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@467 N_OUT7_Mp7@467_d N_OUT6_Mp7@467_g N_VDD_Mp7@467_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@466 N_OUT7_Mp7@466_d N_OUT6_Mp7@466_g N_VDD_Mp7@466_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@465 N_OUT7_Mn7@465_d N_OUT6_Mn7@465_g N_VSS_Mn7@465_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@464 N_OUT7_Mn7@464_d N_OUT6_Mn7@464_g N_VSS_Mn7@464_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@465 N_OUT7_Mp7@465_d N_OUT6_Mp7@465_g N_VDD_Mp7@465_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@464 N_OUT7_Mp7@464_d N_OUT6_Mp7@464_g N_VDD_Mp7@464_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@463 N_OUT7_Mn7@463_d N_OUT6_Mn7@463_g N_VSS_Mn7@463_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@462 N_OUT7_Mn7@462_d N_OUT6_Mn7@462_g N_VSS_Mn7@462_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@463 N_OUT7_Mp7@463_d N_OUT6_Mp7@463_g N_VDD_Mp7@463_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@462 N_OUT7_Mp7@462_d N_OUT6_Mp7@462_g N_VDD_Mp7@462_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@461 N_OUT7_Mn7@461_d N_OUT6_Mn7@461_g N_VSS_Mn7@461_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@460 N_OUT7_Mn7@460_d N_OUT6_Mn7@460_g N_VSS_Mn7@460_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@461 N_OUT7_Mp7@461_d N_OUT6_Mp7@461_g N_VDD_Mp7@461_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@460 N_OUT7_Mp7@460_d N_OUT6_Mp7@460_g N_VDD_Mp7@460_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@459 N_OUT7_Mn7@459_d N_OUT6_Mn7@459_g N_VSS_Mn7@459_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@458 N_OUT7_Mn7@458_d N_OUT6_Mn7@458_g N_VSS_Mn7@458_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@459 N_OUT7_Mp7@459_d N_OUT6_Mp7@459_g N_VDD_Mp7@459_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@458 N_OUT7_Mp7@458_d N_OUT6_Mp7@458_g N_VDD_Mp7@458_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@457 N_OUT7_Mn7@457_d N_OUT6_Mn7@457_g N_VSS_Mn7@457_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@456 N_OUT7_Mn7@456_d N_OUT6_Mn7@456_g N_VSS_Mn7@456_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@457 N_OUT7_Mp7@457_d N_OUT6_Mp7@457_g N_VDD_Mp7@457_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@456 N_OUT7_Mp7@456_d N_OUT6_Mp7@456_g N_VDD_Mp7@456_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@455 N_OUT7_Mn7@455_d N_OUT6_Mn7@455_g N_VSS_Mn7@455_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@454 N_OUT7_Mn7@454_d N_OUT6_Mn7@454_g N_VSS_Mn7@454_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@455 N_OUT7_Mp7@455_d N_OUT6_Mp7@455_g N_VDD_Mp7@455_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@454 N_OUT7_Mp7@454_d N_OUT6_Mp7@454_g N_VDD_Mp7@454_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@453 N_OUT7_Mn7@453_d N_OUT6_Mn7@453_g N_VSS_Mn7@453_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@452 N_OUT7_Mn7@452_d N_OUT6_Mn7@452_g N_VSS_Mn7@452_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@453 N_OUT7_Mp7@453_d N_OUT6_Mp7@453_g N_VDD_Mp7@453_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@452 N_OUT7_Mp7@452_d N_OUT6_Mp7@452_g N_VDD_Mp7@452_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@451 N_OUT7_Mn7@451_d N_OUT6_Mn7@451_g N_VSS_Mn7@451_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@450 N_OUT7_Mn7@450_d N_OUT6_Mn7@450_g N_VSS_Mn7@450_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@451 N_OUT7_Mp7@451_d N_OUT6_Mp7@451_g N_VDD_Mp7@451_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@450 N_OUT7_Mp7@450_d N_OUT6_Mp7@450_g N_VDD_Mp7@450_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@449 N_OUT7_Mn7@449_d N_OUT6_Mn7@449_g N_VSS_Mn7@449_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@448 N_OUT7_Mn7@448_d N_OUT6_Mn7@448_g N_VSS_Mn7@448_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@449 N_OUT7_Mp7@449_d N_OUT6_Mp7@449_g N_VDD_Mp7@449_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@448 N_OUT7_Mp7@448_d N_OUT6_Mp7@448_g N_VDD_Mp7@448_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@447 N_OUT7_Mn7@447_d N_OUT6_Mn7@447_g N_VSS_Mn7@447_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@446 N_OUT7_Mn7@446_d N_OUT6_Mn7@446_g N_VSS_Mn7@446_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@447 N_OUT7_Mp7@447_d N_OUT6_Mp7@447_g N_VDD_Mp7@447_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@446 N_OUT7_Mp7@446_d N_OUT6_Mp7@446_g N_VDD_Mp7@446_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@445 N_OUT7_Mn7@445_d N_OUT6_Mn7@445_g N_VSS_Mn7@445_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@444 N_OUT7_Mn7@444_d N_OUT6_Mn7@444_g N_VSS_Mn7@444_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@445 N_OUT7_Mp7@445_d N_OUT6_Mp7@445_g N_VDD_Mp7@445_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@444 N_OUT7_Mp7@444_d N_OUT6_Mp7@444_g N_VDD_Mp7@444_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@443 N_OUT7_Mn7@443_d N_OUT6_Mn7@443_g N_VSS_Mn7@443_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@442 N_OUT7_Mn7@442_d N_OUT6_Mn7@442_g N_VSS_Mn7@442_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@443 N_OUT7_Mp7@443_d N_OUT6_Mp7@443_g N_VDD_Mp7@443_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@442 N_OUT7_Mp7@442_d N_OUT6_Mp7@442_g N_VDD_Mp7@442_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@441 N_OUT7_Mn7@441_d N_OUT6_Mn7@441_g N_VSS_Mn7@441_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@440 N_OUT7_Mn7@440_d N_OUT6_Mn7@440_g N_VSS_Mn7@440_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@441 N_OUT7_Mp7@441_d N_OUT6_Mp7@441_g N_VDD_Mp7@441_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@440 N_OUT7_Mp7@440_d N_OUT6_Mp7@440_g N_VDD_Mp7@440_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@439 N_OUT7_Mn7@439_d N_OUT6_Mn7@439_g N_VSS_Mn7@439_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@438 N_OUT7_Mn7@438_d N_OUT6_Mn7@438_g N_VSS_Mn7@438_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@439 N_OUT7_Mp7@439_d N_OUT6_Mp7@439_g N_VDD_Mp7@439_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@438 N_OUT7_Mp7@438_d N_OUT6_Mp7@438_g N_VDD_Mp7@438_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@437 N_OUT7_Mn7@437_d N_OUT6_Mn7@437_g N_VSS_Mn7@437_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@436 N_OUT7_Mn7@436_d N_OUT6_Mn7@436_g N_VSS_Mn7@436_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@437 N_OUT7_Mp7@437_d N_OUT6_Mp7@437_g N_VDD_Mp7@437_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@436 N_OUT7_Mp7@436_d N_OUT6_Mp7@436_g N_VDD_Mp7@436_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@435 N_OUT7_Mn7@435_d N_OUT6_Mn7@435_g N_VSS_Mn7@435_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@434 N_OUT7_Mn7@434_d N_OUT6_Mn7@434_g N_VSS_Mn7@434_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@435 N_OUT7_Mp7@435_d N_OUT6_Mp7@435_g N_VDD_Mp7@435_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@434 N_OUT7_Mp7@434_d N_OUT6_Mp7@434_g N_VDD_Mp7@434_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@433 N_OUT7_Mn7@433_d N_OUT6_Mn7@433_g N_VSS_Mn7@433_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@432 N_OUT7_Mn7@432_d N_OUT6_Mn7@432_g N_VSS_Mn7@432_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@433 N_OUT7_Mp7@433_d N_OUT6_Mp7@433_g N_VDD_Mp7@433_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@432 N_OUT7_Mp7@432_d N_OUT6_Mp7@432_g N_VDD_Mp7@432_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@431 N_OUT7_Mn7@431_d N_OUT6_Mn7@431_g N_VSS_Mn7@431_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@430 N_OUT7_Mn7@430_d N_OUT6_Mn7@430_g N_VSS_Mn7@430_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@431 N_OUT7_Mp7@431_d N_OUT6_Mp7@431_g N_VDD_Mp7@431_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@430 N_OUT7_Mp7@430_d N_OUT6_Mp7@430_g N_VDD_Mp7@430_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@429 N_OUT7_Mn7@429_d N_OUT6_Mn7@429_g N_VSS_Mn7@429_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@428 N_OUT7_Mn7@428_d N_OUT6_Mn7@428_g N_VSS_Mn7@428_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@429 N_OUT7_Mp7@429_d N_OUT6_Mp7@429_g N_VDD_Mp7@429_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@428 N_OUT7_Mp7@428_d N_OUT6_Mp7@428_g N_VDD_Mp7@428_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@427 N_OUT7_Mn7@427_d N_OUT6_Mn7@427_g N_VSS_Mn7@427_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@426 N_OUT7_Mn7@426_d N_OUT6_Mn7@426_g N_VSS_Mn7@426_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@427 N_OUT7_Mp7@427_d N_OUT6_Mp7@427_g N_VDD_Mp7@427_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@426 N_OUT7_Mp7@426_d N_OUT6_Mp7@426_g N_VDD_Mp7@426_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@425 N_OUT7_Mn7@425_d N_OUT6_Mn7@425_g N_VSS_Mn7@425_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@424 N_OUT7_Mn7@424_d N_OUT6_Mn7@424_g N_VSS_Mn7@424_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@425 N_OUT7_Mp7@425_d N_OUT6_Mp7@425_g N_VDD_Mp7@425_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@424 N_OUT7_Mp7@424_d N_OUT6_Mp7@424_g N_VDD_Mp7@424_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@423 N_OUT7_Mn7@423_d N_OUT6_Mn7@423_g N_VSS_Mn7@423_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@422 N_OUT7_Mn7@422_d N_OUT6_Mn7@422_g N_VSS_Mn7@422_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@423 N_OUT7_Mp7@423_d N_OUT6_Mp7@423_g N_VDD_Mp7@423_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@422 N_OUT7_Mp7@422_d N_OUT6_Mp7@422_g N_VDD_Mp7@422_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@421 N_OUT7_Mn7@421_d N_OUT6_Mn7@421_g N_VSS_Mn7@421_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@420 N_OUT7_Mn7@420_d N_OUT6_Mn7@420_g N_VSS_Mn7@420_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@421 N_OUT7_Mp7@421_d N_OUT6_Mp7@421_g N_VDD_Mp7@421_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@420 N_OUT7_Mp7@420_d N_OUT6_Mp7@420_g N_VDD_Mp7@420_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@419 N_OUT7_Mn7@419_d N_OUT6_Mn7@419_g N_VSS_Mn7@419_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@418 N_OUT7_Mn7@418_d N_OUT6_Mn7@418_g N_VSS_Mn7@418_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@419 N_OUT7_Mp7@419_d N_OUT6_Mp7@419_g N_VDD_Mp7@419_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@418 N_OUT7_Mp7@418_d N_OUT6_Mp7@418_g N_VDD_Mp7@418_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@417 N_OUT7_Mn7@417_d N_OUT6_Mn7@417_g N_VSS_Mn7@417_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@416 N_OUT7_Mn7@416_d N_OUT6_Mn7@416_g N_VSS_Mn7@416_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@417 N_OUT7_Mp7@417_d N_OUT6_Mp7@417_g N_VDD_Mp7@417_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@416 N_OUT7_Mp7@416_d N_OUT6_Mp7@416_g N_VDD_Mp7@416_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@415 N_OUT7_Mn7@415_d N_OUT6_Mn7@415_g N_VSS_Mn7@415_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@414 N_OUT7_Mn7@414_d N_OUT6_Mn7@414_g N_VSS_Mn7@414_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@415 N_OUT7_Mp7@415_d N_OUT6_Mp7@415_g N_VDD_Mp7@415_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@414 N_OUT7_Mp7@414_d N_OUT6_Mp7@414_g N_VDD_Mp7@414_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@413 N_OUT7_Mn7@413_d N_OUT6_Mn7@413_g N_VSS_Mn7@413_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@412 N_OUT7_Mn7@412_d N_OUT6_Mn7@412_g N_VSS_Mn7@412_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@413 N_OUT7_Mp7@413_d N_OUT6_Mp7@413_g N_VDD_Mp7@413_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@412 N_OUT7_Mp7@412_d N_OUT6_Mp7@412_g N_VDD_Mp7@412_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@411 N_OUT7_Mn7@411_d N_OUT6_Mn7@411_g N_VSS_Mn7@411_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@410 N_OUT7_Mn7@410_d N_OUT6_Mn7@410_g N_VSS_Mn7@410_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@411 N_OUT7_Mp7@411_d N_OUT6_Mp7@411_g N_VDD_Mp7@411_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@410 N_OUT7_Mp7@410_d N_OUT6_Mp7@410_g N_VDD_Mp7@410_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@409 N_OUT7_Mn7@409_d N_OUT6_Mn7@409_g N_VSS_Mn7@409_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@408 N_OUT7_Mn7@408_d N_OUT6_Mn7@408_g N_VSS_Mn7@408_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@409 N_OUT7_Mp7@409_d N_OUT6_Mp7@409_g N_VDD_Mp7@409_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@408 N_OUT7_Mp7@408_d N_OUT6_Mp7@408_g N_VDD_Mp7@408_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@407 N_OUT7_Mn7@407_d N_OUT6_Mn7@407_g N_VSS_Mn7@407_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@406 N_OUT7_Mn7@406_d N_OUT6_Mn7@406_g N_VSS_Mn7@406_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@407 N_OUT7_Mp7@407_d N_OUT6_Mp7@407_g N_VDD_Mp7@407_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@406 N_OUT7_Mp7@406_d N_OUT6_Mp7@406_g N_VDD_Mp7@406_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@405 N_OUT7_Mn7@405_d N_OUT6_Mn7@405_g N_VSS_Mn7@405_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@404 N_OUT7_Mn7@404_d N_OUT6_Mn7@404_g N_VSS_Mn7@404_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@405 N_OUT7_Mp7@405_d N_OUT6_Mp7@405_g N_VDD_Mp7@405_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@404 N_OUT7_Mp7@404_d N_OUT6_Mp7@404_g N_VDD_Mp7@404_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@403 N_OUT7_Mn7@403_d N_OUT6_Mn7@403_g N_VSS_Mn7@403_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@402 N_OUT7_Mn7@402_d N_OUT6_Mn7@402_g N_VSS_Mn7@402_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@403 N_OUT7_Mp7@403_d N_OUT6_Mp7@403_g N_VDD_Mp7@403_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@402 N_OUT7_Mp7@402_d N_OUT6_Mp7@402_g N_VDD_Mp7@402_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@401 N_OUT7_Mn7@401_d N_OUT6_Mn7@401_g N_VSS_Mn7@401_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@400 N_OUT7_Mn7@400_d N_OUT6_Mn7@400_g N_VSS_Mn7@400_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@401 N_OUT7_Mp7@401_d N_OUT6_Mp7@401_g N_VDD_Mp7@401_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@400 N_OUT7_Mp7@400_d N_OUT6_Mp7@400_g N_VDD_Mp7@400_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@399 N_OUT7_Mn7@399_d N_OUT6_Mn7@399_g N_VSS_Mn7@399_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@398 N_OUT7_Mn7@398_d N_OUT6_Mn7@398_g N_VSS_Mn7@398_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@399 N_OUT7_Mp7@399_d N_OUT6_Mp7@399_g N_VDD_Mp7@399_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@398 N_OUT7_Mp7@398_d N_OUT6_Mp7@398_g N_VDD_Mp7@398_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@397 N_OUT7_Mn7@397_d N_OUT6_Mn7@397_g N_VSS_Mn7@397_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@396 N_OUT7_Mn7@396_d N_OUT6_Mn7@396_g N_VSS_Mn7@396_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@397 N_OUT7_Mp7@397_d N_OUT6_Mp7@397_g N_VDD_Mp7@397_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@396 N_OUT7_Mp7@396_d N_OUT6_Mp7@396_g N_VDD_Mp7@396_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@395 N_OUT7_Mn7@395_d N_OUT6_Mn7@395_g N_VSS_Mn7@395_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@394 N_OUT7_Mn7@394_d N_OUT6_Mn7@394_g N_VSS_Mn7@394_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@395 N_OUT7_Mp7@395_d N_OUT6_Mp7@395_g N_VDD_Mp7@395_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@394 N_OUT7_Mp7@394_d N_OUT6_Mp7@394_g N_VDD_Mp7@394_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@393 N_OUT7_Mn7@393_d N_OUT6_Mn7@393_g N_VSS_Mn7@393_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@392 N_OUT7_Mn7@392_d N_OUT6_Mn7@392_g N_VSS_Mn7@392_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@393 N_OUT7_Mp7@393_d N_OUT6_Mp7@393_g N_VDD_Mp7@393_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@392 N_OUT7_Mp7@392_d N_OUT6_Mp7@392_g N_VDD_Mp7@392_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@391 N_OUT7_Mn7@391_d N_OUT6_Mn7@391_g N_VSS_Mn7@391_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@390 N_OUT7_Mn7@390_d N_OUT6_Mn7@390_g N_VSS_Mn7@390_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@391 N_OUT7_Mp7@391_d N_OUT6_Mp7@391_g N_VDD_Mp7@391_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@390 N_OUT7_Mp7@390_d N_OUT6_Mp7@390_g N_VDD_Mp7@390_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@389 N_OUT7_Mn7@389_d N_OUT6_Mn7@389_g N_VSS_Mn7@389_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@388 N_OUT7_Mn7@388_d N_OUT6_Mn7@388_g N_VSS_Mn7@388_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@389 N_OUT7_Mp7@389_d N_OUT6_Mp7@389_g N_VDD_Mp7@389_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@388 N_OUT7_Mp7@388_d N_OUT6_Mp7@388_g N_VDD_Mp7@388_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@387 N_OUT7_Mn7@387_d N_OUT6_Mn7@387_g N_VSS_Mn7@387_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@386 N_OUT7_Mn7@386_d N_OUT6_Mn7@386_g N_VSS_Mn7@386_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@387 N_OUT7_Mp7@387_d N_OUT6_Mp7@387_g N_VDD_Mp7@387_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@386 N_OUT7_Mp7@386_d N_OUT6_Mp7@386_g N_VDD_Mp7@386_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@385 N_OUT7_Mn7@385_d N_OUT6_Mn7@385_g N_VSS_Mn7@385_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@384 N_OUT7_Mn7@384_d N_OUT6_Mn7@384_g N_VSS_Mn7@384_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@385 N_OUT7_Mp7@385_d N_OUT6_Mp7@385_g N_VDD_Mp7@385_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@384 N_OUT7_Mp7@384_d N_OUT6_Mp7@384_g N_VDD_Mp7@384_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@383 N_OUT7_Mn7@383_d N_OUT6_Mn7@383_g N_VSS_Mn7@383_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@382 N_OUT7_Mn7@382_d N_OUT6_Mn7@382_g N_VSS_Mn7@382_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@383 N_OUT7_Mp7@383_d N_OUT6_Mp7@383_g N_VDD_Mp7@383_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@382 N_OUT7_Mp7@382_d N_OUT6_Mp7@382_g N_VDD_Mp7@382_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@381 N_OUT7_Mn7@381_d N_OUT6_Mn7@381_g N_VSS_Mn7@381_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@380 N_OUT7_Mn7@380_d N_OUT6_Mn7@380_g N_VSS_Mn7@380_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@381 N_OUT7_Mp7@381_d N_OUT6_Mp7@381_g N_VDD_Mp7@381_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@380 N_OUT7_Mp7@380_d N_OUT6_Mp7@380_g N_VDD_Mp7@380_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@379 N_OUT7_Mn7@379_d N_OUT6_Mn7@379_g N_VSS_Mn7@379_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@378 N_OUT7_Mn7@378_d N_OUT6_Mn7@378_g N_VSS_Mn7@378_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@379 N_OUT7_Mp7@379_d N_OUT6_Mp7@379_g N_VDD_Mp7@379_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@378 N_OUT7_Mp7@378_d N_OUT6_Mp7@378_g N_VDD_Mp7@378_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@377 N_OUT7_Mn7@377_d N_OUT6_Mn7@377_g N_VSS_Mn7@377_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@376 N_OUT7_Mn7@376_d N_OUT6_Mn7@376_g N_VSS_Mn7@376_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@377 N_OUT7_Mp7@377_d N_OUT6_Mp7@377_g N_VDD_Mp7@377_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@376 N_OUT7_Mp7@376_d N_OUT6_Mp7@376_g N_VDD_Mp7@376_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@375 N_OUT7_Mn7@375_d N_OUT6_Mn7@375_g N_VSS_Mn7@375_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@374 N_OUT7_Mn7@374_d N_OUT6_Mn7@374_g N_VSS_Mn7@374_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@375 N_OUT7_Mp7@375_d N_OUT6_Mp7@375_g N_VDD_Mp7@375_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@374 N_OUT7_Mp7@374_d N_OUT6_Mp7@374_g N_VDD_Mp7@374_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@373 N_OUT7_Mn7@373_d N_OUT6_Mn7@373_g N_VSS_Mn7@373_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@372 N_OUT7_Mn7@372_d N_OUT6_Mn7@372_g N_VSS_Mn7@372_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@373 N_OUT7_Mp7@373_d N_OUT6_Mp7@373_g N_VDD_Mp7@373_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@372 N_OUT7_Mp7@372_d N_OUT6_Mp7@372_g N_VDD_Mp7@372_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@371 N_OUT7_Mn7@371_d N_OUT6_Mn7@371_g N_VSS_Mn7@371_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@370 N_OUT7_Mn7@370_d N_OUT6_Mn7@370_g N_VSS_Mn7@370_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@371 N_OUT7_Mp7@371_d N_OUT6_Mp7@371_g N_VDD_Mp7@371_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@370 N_OUT7_Mp7@370_d N_OUT6_Mp7@370_g N_VDD_Mp7@370_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@369 N_OUT7_Mn7@369_d N_OUT6_Mn7@369_g N_VSS_Mn7@369_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@368 N_OUT7_Mn7@368_d N_OUT6_Mn7@368_g N_VSS_Mn7@368_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@369 N_OUT7_Mp7@369_d N_OUT6_Mp7@369_g N_VDD_Mp7@369_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@368 N_OUT7_Mp7@368_d N_OUT6_Mp7@368_g N_VDD_Mp7@368_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@367 N_OUT7_Mn7@367_d N_OUT6_Mn7@367_g N_VSS_Mn7@367_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@366 N_OUT7_Mn7@366_d N_OUT6_Mn7@366_g N_VSS_Mn7@366_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@367 N_OUT7_Mp7@367_d N_OUT6_Mp7@367_g N_VDD_Mp7@367_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@366 N_OUT7_Mp7@366_d N_OUT6_Mp7@366_g N_VDD_Mp7@366_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@365 N_OUT7_Mn7@365_d N_OUT6_Mn7@365_g N_VSS_Mn7@365_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@364 N_OUT7_Mn7@364_d N_OUT6_Mn7@364_g N_VSS_Mn7@364_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@365 N_OUT7_Mp7@365_d N_OUT6_Mp7@365_g N_VDD_Mp7@365_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@364 N_OUT7_Mp7@364_d N_OUT6_Mp7@364_g N_VDD_Mp7@364_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@363 N_OUT7_Mn7@363_d N_OUT6_Mn7@363_g N_VSS_Mn7@363_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@362 N_OUT7_Mn7@362_d N_OUT6_Mn7@362_g N_VSS_Mn7@362_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@363 N_OUT7_Mp7@363_d N_OUT6_Mp7@363_g N_VDD_Mp7@363_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@362 N_OUT7_Mp7@362_d N_OUT6_Mp7@362_g N_VDD_Mp7@362_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@361 N_OUT7_Mn7@361_d N_OUT6_Mn7@361_g N_VSS_Mn7@361_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@360 N_OUT7_Mn7@360_d N_OUT6_Mn7@360_g N_VSS_Mn7@360_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@361 N_OUT7_Mp7@361_d N_OUT6_Mp7@361_g N_VDD_Mp7@361_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@360 N_OUT7_Mp7@360_d N_OUT6_Mp7@360_g N_VDD_Mp7@360_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@359 N_OUT7_Mn7@359_d N_OUT6_Mn7@359_g N_VSS_Mn7@359_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@358 N_OUT7_Mn7@358_d N_OUT6_Mn7@358_g N_VSS_Mn7@358_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@359 N_OUT7_Mp7@359_d N_OUT6_Mp7@359_g N_VDD_Mp7@359_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@358 N_OUT7_Mp7@358_d N_OUT6_Mp7@358_g N_VDD_Mp7@358_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@357 N_OUT7_Mn7@357_d N_OUT6_Mn7@357_g N_VSS_Mn7@357_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@356 N_OUT7_Mn7@356_d N_OUT6_Mn7@356_g N_VSS_Mn7@356_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@357 N_OUT7_Mp7@357_d N_OUT6_Mp7@357_g N_VDD_Mp7@357_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@356 N_OUT7_Mp7@356_d N_OUT6_Mp7@356_g N_VDD_Mp7@356_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@355 N_OUT7_Mn7@355_d N_OUT6_Mn7@355_g N_VSS_Mn7@355_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@354 N_OUT7_Mn7@354_d N_OUT6_Mn7@354_g N_VSS_Mn7@354_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@355 N_OUT7_Mp7@355_d N_OUT6_Mp7@355_g N_VDD_Mp7@355_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@354 N_OUT7_Mp7@354_d N_OUT6_Mp7@354_g N_VDD_Mp7@354_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@353 N_OUT7_Mn7@353_d N_OUT6_Mn7@353_g N_VSS_Mn7@353_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@352 N_OUT7_Mn7@352_d N_OUT6_Mn7@352_g N_VSS_Mn7@352_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@353 N_OUT7_Mp7@353_d N_OUT6_Mp7@353_g N_VDD_Mp7@353_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@352 N_OUT7_Mp7@352_d N_OUT6_Mp7@352_g N_VDD_Mp7@352_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@351 N_OUT7_Mn7@351_d N_OUT6_Mn7@351_g N_VSS_Mn7@351_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@350 N_OUT7_Mn7@350_d N_OUT6_Mn7@350_g N_VSS_Mn7@350_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@351 N_OUT7_Mp7@351_d N_OUT6_Mp7@351_g N_VDD_Mp7@351_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@350 N_OUT7_Mp7@350_d N_OUT6_Mp7@350_g N_VDD_Mp7@350_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@349 N_OUT7_Mn7@349_d N_OUT6_Mn7@349_g N_VSS_Mn7@349_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@348 N_OUT7_Mn7@348_d N_OUT6_Mn7@348_g N_VSS_Mn7@348_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@349 N_OUT7_Mp7@349_d N_OUT6_Mp7@349_g N_VDD_Mp7@349_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@348 N_OUT7_Mp7@348_d N_OUT6_Mp7@348_g N_VDD_Mp7@348_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@347 N_OUT7_Mn7@347_d N_OUT6_Mn7@347_g N_VSS_Mn7@347_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@346 N_OUT7_Mn7@346_d N_OUT6_Mn7@346_g N_VSS_Mn7@346_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@347 N_OUT7_Mp7@347_d N_OUT6_Mp7@347_g N_VDD_Mp7@347_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@346 N_OUT7_Mp7@346_d N_OUT6_Mp7@346_g N_VDD_Mp7@346_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@345 N_OUT7_Mn7@345_d N_OUT6_Mn7@345_g N_VSS_Mn7@345_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@344 N_OUT7_Mn7@344_d N_OUT6_Mn7@344_g N_VSS_Mn7@344_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@345 N_OUT7_Mp7@345_d N_OUT6_Mp7@345_g N_VDD_Mp7@345_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@344 N_OUT7_Mp7@344_d N_OUT6_Mp7@344_g N_VDD_Mp7@344_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@343 N_OUT7_Mn7@343_d N_OUT6_Mn7@343_g N_VSS_Mn7@343_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@342 N_OUT7_Mn7@342_d N_OUT6_Mn7@342_g N_VSS_Mn7@342_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@343 N_OUT7_Mp7@343_d N_OUT6_Mp7@343_g N_VDD_Mp7@343_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@342 N_OUT7_Mp7@342_d N_OUT6_Mp7@342_g N_VDD_Mp7@342_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@341 N_OUT7_Mn7@341_d N_OUT6_Mn7@341_g N_VSS_Mn7@341_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@340 N_OUT7_Mn7@340_d N_OUT6_Mn7@340_g N_VSS_Mn7@340_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@341 N_OUT7_Mp7@341_d N_OUT6_Mp7@341_g N_VDD_Mp7@341_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@340 N_OUT7_Mp7@340_d N_OUT6_Mp7@340_g N_VDD_Mp7@340_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@339 N_OUT7_Mn7@339_d N_OUT6_Mn7@339_g N_VSS_Mn7@339_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@338 N_OUT7_Mn7@338_d N_OUT6_Mn7@338_g N_VSS_Mn7@338_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@339 N_OUT7_Mp7@339_d N_OUT6_Mp7@339_g N_VDD_Mp7@339_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@338 N_OUT7_Mp7@338_d N_OUT6_Mp7@338_g N_VDD_Mp7@338_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@337 N_OUT7_Mn7@337_d N_OUT6_Mn7@337_g N_VSS_Mn7@337_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@336 N_OUT7_Mn7@336_d N_OUT6_Mn7@336_g N_VSS_Mn7@336_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@337 N_OUT7_Mp7@337_d N_OUT6_Mp7@337_g N_VDD_Mp7@337_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@336 N_OUT7_Mp7@336_d N_OUT6_Mp7@336_g N_VDD_Mp7@336_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@335 N_OUT7_Mn7@335_d N_OUT6_Mn7@335_g N_VSS_Mn7@335_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@334 N_OUT7_Mn7@334_d N_OUT6_Mn7@334_g N_VSS_Mn7@334_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@335 N_OUT7_Mp7@335_d N_OUT6_Mp7@335_g N_VDD_Mp7@335_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@334 N_OUT7_Mp7@334_d N_OUT6_Mp7@334_g N_VDD_Mp7@334_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@333 N_OUT7_Mn7@333_d N_OUT6_Mn7@333_g N_VSS_Mn7@333_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@332 N_OUT7_Mn7@332_d N_OUT6_Mn7@332_g N_VSS_Mn7@332_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@333 N_OUT7_Mp7@333_d N_OUT6_Mp7@333_g N_VDD_Mp7@333_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@332 N_OUT7_Mp7@332_d N_OUT6_Mp7@332_g N_VDD_Mp7@332_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@331 N_OUT7_Mn7@331_d N_OUT6_Mn7@331_g N_VSS_Mn7@331_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@330 N_OUT7_Mn7@330_d N_OUT6_Mn7@330_g N_VSS_Mn7@330_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@331 N_OUT7_Mp7@331_d N_OUT6_Mp7@331_g N_VDD_Mp7@331_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@330 N_OUT7_Mp7@330_d N_OUT6_Mp7@330_g N_VDD_Mp7@330_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@329 N_OUT7_Mn7@329_d N_OUT6_Mn7@329_g N_VSS_Mn7@329_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@328 N_OUT7_Mn7@328_d N_OUT6_Mn7@328_g N_VSS_Mn7@328_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@329 N_OUT7_Mp7@329_d N_OUT6_Mp7@329_g N_VDD_Mp7@329_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@328 N_OUT7_Mp7@328_d N_OUT6_Mp7@328_g N_VDD_Mp7@328_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@327 N_OUT7_Mn7@327_d N_OUT6_Mn7@327_g N_VSS_Mn7@327_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@326 N_OUT7_Mn7@326_d N_OUT6_Mn7@326_g N_VSS_Mn7@326_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@327 N_OUT7_Mp7@327_d N_OUT6_Mp7@327_g N_VDD_Mp7@327_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@326 N_OUT7_Mp7@326_d N_OUT6_Mp7@326_g N_VDD_Mp7@326_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@325 N_OUT7_Mn7@325_d N_OUT6_Mn7@325_g N_VSS_Mn7@325_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@324 N_OUT7_Mn7@324_d N_OUT6_Mn7@324_g N_VSS_Mn7@324_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@325 N_OUT7_Mp7@325_d N_OUT6_Mp7@325_g N_VDD_Mp7@325_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@324 N_OUT7_Mp7@324_d N_OUT6_Mp7@324_g N_VDD_Mp7@324_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@323 N_OUT7_Mn7@323_d N_OUT6_Mn7@323_g N_VSS_Mn7@323_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@322 N_OUT7_Mn7@322_d N_OUT6_Mn7@322_g N_VSS_Mn7@322_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@323 N_OUT7_Mp7@323_d N_OUT6_Mp7@323_g N_VDD_Mp7@323_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@322 N_OUT7_Mp7@322_d N_OUT6_Mp7@322_g N_VDD_Mp7@322_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@321 N_OUT7_Mn7@321_d N_OUT6_Mn7@321_g N_VSS_Mn7@321_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@320 N_OUT7_Mn7@320_d N_OUT6_Mn7@320_g N_VSS_Mn7@320_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@321 N_OUT7_Mp7@321_d N_OUT6_Mp7@321_g N_VDD_Mp7@321_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@320 N_OUT7_Mp7@320_d N_OUT6_Mp7@320_g N_VDD_Mp7@320_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@319 N_OUT7_Mn7@319_d N_OUT6_Mn7@319_g N_VSS_Mn7@319_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@318 N_OUT7_Mn7@318_d N_OUT6_Mn7@318_g N_VSS_Mn7@318_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@319 N_OUT7_Mp7@319_d N_OUT6_Mp7@319_g N_VDD_Mp7@319_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@318 N_OUT7_Mp7@318_d N_OUT6_Mp7@318_g N_VDD_Mp7@318_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@317 N_OUT7_Mn7@317_d N_OUT6_Mn7@317_g N_VSS_Mn7@317_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@316 N_OUT7_Mn7@316_d N_OUT6_Mn7@316_g N_VSS_Mn7@316_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@317 N_OUT7_Mp7@317_d N_OUT6_Mp7@317_g N_VDD_Mp7@317_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@316 N_OUT7_Mp7@316_d N_OUT6_Mp7@316_g N_VDD_Mp7@316_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@315 N_OUT7_Mn7@315_d N_OUT6_Mn7@315_g N_VSS_Mn7@315_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@314 N_OUT7_Mn7@314_d N_OUT6_Mn7@314_g N_VSS_Mn7@314_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@315 N_OUT7_Mp7@315_d N_OUT6_Mp7@315_g N_VDD_Mp7@315_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@314 N_OUT7_Mp7@314_d N_OUT6_Mp7@314_g N_VDD_Mp7@314_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@313 N_OUT7_Mn7@313_d N_OUT6_Mn7@313_g N_VSS_Mn7@313_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@312 N_OUT7_Mn7@312_d N_OUT6_Mn7@312_g N_VSS_Mn7@312_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@313 N_OUT7_Mp7@313_d N_OUT6_Mp7@313_g N_VDD_Mp7@313_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@312 N_OUT7_Mp7@312_d N_OUT6_Mp7@312_g N_VDD_Mp7@312_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@311 N_OUT7_Mn7@311_d N_OUT6_Mn7@311_g N_VSS_Mn7@311_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@310 N_OUT7_Mn7@310_d N_OUT6_Mn7@310_g N_VSS_Mn7@310_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@311 N_OUT7_Mp7@311_d N_OUT6_Mp7@311_g N_VDD_Mp7@311_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@310 N_OUT7_Mp7@310_d N_OUT6_Mp7@310_g N_VDD_Mp7@310_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@309 N_OUT7_Mn7@309_d N_OUT6_Mn7@309_g N_VSS_Mn7@309_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@308 N_OUT7_Mn7@308_d N_OUT6_Mn7@308_g N_VSS_Mn7@308_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@309 N_OUT7_Mp7@309_d N_OUT6_Mp7@309_g N_VDD_Mp7@309_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@308 N_OUT7_Mp7@308_d N_OUT6_Mp7@308_g N_VDD_Mp7@308_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@307 N_OUT7_Mn7@307_d N_OUT6_Mn7@307_g N_VSS_Mn7@307_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@306 N_OUT7_Mn7@306_d N_OUT6_Mn7@306_g N_VSS_Mn7@306_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@307 N_OUT7_Mp7@307_d N_OUT6_Mp7@307_g N_VDD_Mp7@307_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@306 N_OUT7_Mp7@306_d N_OUT6_Mp7@306_g N_VDD_Mp7@306_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@305 N_OUT7_Mn7@305_d N_OUT6_Mn7@305_g N_VSS_Mn7@305_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@304 N_OUT7_Mn7@304_d N_OUT6_Mn7@304_g N_VSS_Mn7@304_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@305 N_OUT7_Mp7@305_d N_OUT6_Mp7@305_g N_VDD_Mp7@305_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@304 N_OUT7_Mp7@304_d N_OUT6_Mp7@304_g N_VDD_Mp7@304_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@303 N_OUT7_Mn7@303_d N_OUT6_Mn7@303_g N_VSS_Mn7@303_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@302 N_OUT7_Mn7@302_d N_OUT6_Mn7@302_g N_VSS_Mn7@302_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@303 N_OUT7_Mp7@303_d N_OUT6_Mp7@303_g N_VDD_Mp7@303_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@302 N_OUT7_Mp7@302_d N_OUT6_Mp7@302_g N_VDD_Mp7@302_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@301 N_OUT7_Mn7@301_d N_OUT6_Mn7@301_g N_VSS_Mn7@301_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@300 N_OUT7_Mn7@300_d N_OUT6_Mn7@300_g N_VSS_Mn7@300_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@301 N_OUT7_Mp7@301_d N_OUT6_Mp7@301_g N_VDD_Mp7@301_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@300 N_OUT7_Mp7@300_d N_OUT6_Mp7@300_g N_VDD_Mp7@300_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@299 N_OUT7_Mn7@299_d N_OUT6_Mn7@299_g N_VSS_Mn7@299_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@298 N_OUT7_Mn7@298_d N_OUT6_Mn7@298_g N_VSS_Mn7@298_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@299 N_OUT7_Mp7@299_d N_OUT6_Mp7@299_g N_VDD_Mp7@299_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@298 N_OUT7_Mp7@298_d N_OUT6_Mp7@298_g N_VDD_Mp7@298_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@297 N_OUT7_Mn7@297_d N_OUT6_Mn7@297_g N_VSS_Mn7@297_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@296 N_OUT7_Mn7@296_d N_OUT6_Mn7@296_g N_VSS_Mn7@296_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@297 N_OUT7_Mp7@297_d N_OUT6_Mp7@297_g N_VDD_Mp7@297_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@296 N_OUT7_Mp7@296_d N_OUT6_Mp7@296_g N_VDD_Mp7@296_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@295 N_OUT7_Mn7@295_d N_OUT6_Mn7@295_g N_VSS_Mn7@295_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@294 N_OUT7_Mn7@294_d N_OUT6_Mn7@294_g N_VSS_Mn7@294_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@295 N_OUT7_Mp7@295_d N_OUT6_Mp7@295_g N_VDD_Mp7@295_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@294 N_OUT7_Mp7@294_d N_OUT6_Mp7@294_g N_VDD_Mp7@294_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@293 N_OUT7_Mn7@293_d N_OUT6_Mn7@293_g N_VSS_Mn7@293_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@292 N_OUT7_Mn7@292_d N_OUT6_Mn7@292_g N_VSS_Mn7@292_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@293 N_OUT7_Mp7@293_d N_OUT6_Mp7@293_g N_VDD_Mp7@293_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@292 N_OUT7_Mp7@292_d N_OUT6_Mp7@292_g N_VDD_Mp7@292_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@291 N_OUT7_Mn7@291_d N_OUT6_Mn7@291_g N_VSS_Mn7@291_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@290 N_OUT7_Mn7@290_d N_OUT6_Mn7@290_g N_VSS_Mn7@290_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@291 N_OUT7_Mp7@291_d N_OUT6_Mp7@291_g N_VDD_Mp7@291_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@290 N_OUT7_Mp7@290_d N_OUT6_Mp7@290_g N_VDD_Mp7@290_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@289 N_OUT7_Mn7@289_d N_OUT6_Mn7@289_g N_VSS_Mn7@289_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@288 N_OUT7_Mn7@288_d N_OUT6_Mn7@288_g N_VSS_Mn7@288_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@289 N_OUT7_Mp7@289_d N_OUT6_Mp7@289_g N_VDD_Mp7@289_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@288 N_OUT7_Mp7@288_d N_OUT6_Mp7@288_g N_VDD_Mp7@288_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@287 N_OUT7_Mn7@287_d N_OUT6_Mn7@287_g N_VSS_Mn7@287_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@286 N_OUT7_Mn7@286_d N_OUT6_Mn7@286_g N_VSS_Mn7@286_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@287 N_OUT7_Mp7@287_d N_OUT6_Mp7@287_g N_VDD_Mp7@287_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@286 N_OUT7_Mp7@286_d N_OUT6_Mp7@286_g N_VDD_Mp7@286_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@285 N_OUT7_Mn7@285_d N_OUT6_Mn7@285_g N_VSS_Mn7@285_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@284 N_OUT7_Mn7@284_d N_OUT6_Mn7@284_g N_VSS_Mn7@284_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@285 N_OUT7_Mp7@285_d N_OUT6_Mp7@285_g N_VDD_Mp7@285_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@284 N_OUT7_Mp7@284_d N_OUT6_Mp7@284_g N_VDD_Mp7@284_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@283 N_OUT7_Mn7@283_d N_OUT6_Mn7@283_g N_VSS_Mn7@283_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@282 N_OUT7_Mn7@282_d N_OUT6_Mn7@282_g N_VSS_Mn7@282_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@283 N_OUT7_Mp7@283_d N_OUT6_Mp7@283_g N_VDD_Mp7@283_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@282 N_OUT7_Mp7@282_d N_OUT6_Mp7@282_g N_VDD_Mp7@282_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@281 N_OUT7_Mn7@281_d N_OUT6_Mn7@281_g N_VSS_Mn7@281_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@280 N_OUT7_Mn7@280_d N_OUT6_Mn7@280_g N_VSS_Mn7@280_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@281 N_OUT7_Mp7@281_d N_OUT6_Mp7@281_g N_VDD_Mp7@281_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@280 N_OUT7_Mp7@280_d N_OUT6_Mp7@280_g N_VDD_Mp7@280_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@279 N_OUT7_Mn7@279_d N_OUT6_Mn7@279_g N_VSS_Mn7@279_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@278 N_OUT7_Mn7@278_d N_OUT6_Mn7@278_g N_VSS_Mn7@278_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@279 N_OUT7_Mp7@279_d N_OUT6_Mp7@279_g N_VDD_Mp7@279_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@278 N_OUT7_Mp7@278_d N_OUT6_Mp7@278_g N_VDD_Mp7@278_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@277 N_OUT7_Mn7@277_d N_OUT6_Mn7@277_g N_VSS_Mn7@277_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@276 N_OUT7_Mn7@276_d N_OUT6_Mn7@276_g N_VSS_Mn7@276_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@277 N_OUT7_Mp7@277_d N_OUT6_Mp7@277_g N_VDD_Mp7@277_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@276 N_OUT7_Mp7@276_d N_OUT6_Mp7@276_g N_VDD_Mp7@276_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@275 N_OUT7_Mn7@275_d N_OUT6_Mn7@275_g N_VSS_Mn7@275_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@274 N_OUT7_Mn7@274_d N_OUT6_Mn7@274_g N_VSS_Mn7@274_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@275 N_OUT7_Mp7@275_d N_OUT6_Mp7@275_g N_VDD_Mp7@275_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@274 N_OUT7_Mp7@274_d N_OUT6_Mp7@274_g N_VDD_Mp7@274_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@273 N_OUT7_Mn7@273_d N_OUT6_Mn7@273_g N_VSS_Mn7@273_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@272 N_OUT7_Mn7@272_d N_OUT6_Mn7@272_g N_VSS_Mn7@272_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@273 N_OUT7_Mp7@273_d N_OUT6_Mp7@273_g N_VDD_Mp7@273_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@272 N_OUT7_Mp7@272_d N_OUT6_Mp7@272_g N_VDD_Mp7@272_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@271 N_OUT7_Mn7@271_d N_OUT6_Mn7@271_g N_VSS_Mn7@271_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@270 N_OUT7_Mn7@270_d N_OUT6_Mn7@270_g N_VSS_Mn7@270_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@271 N_OUT7_Mp7@271_d N_OUT6_Mp7@271_g N_VDD_Mp7@271_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@270 N_OUT7_Mp7@270_d N_OUT6_Mp7@270_g N_VDD_Mp7@270_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@269 N_OUT7_Mn7@269_d N_OUT6_Mn7@269_g N_VSS_Mn7@269_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@268 N_OUT7_Mn7@268_d N_OUT6_Mn7@268_g N_VSS_Mn7@268_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@269 N_OUT7_Mp7@269_d N_OUT6_Mp7@269_g N_VDD_Mp7@269_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@268 N_OUT7_Mp7@268_d N_OUT6_Mp7@268_g N_VDD_Mp7@268_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@267 N_OUT7_Mn7@267_d N_OUT6_Mn7@267_g N_VSS_Mn7@267_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@266 N_OUT7_Mn7@266_d N_OUT6_Mn7@266_g N_VSS_Mn7@266_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@267 N_OUT7_Mp7@267_d N_OUT6_Mp7@267_g N_VDD_Mp7@267_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@266 N_OUT7_Mp7@266_d N_OUT6_Mp7@266_g N_VDD_Mp7@266_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@265 N_OUT7_Mn7@265_d N_OUT6_Mn7@265_g N_VSS_Mn7@265_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@264 N_OUT7_Mn7@264_d N_OUT6_Mn7@264_g N_VSS_Mn7@264_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@265 N_OUT7_Mp7@265_d N_OUT6_Mp7@265_g N_VDD_Mp7@265_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@264 N_OUT7_Mp7@264_d N_OUT6_Mp7@264_g N_VDD_Mp7@264_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@263 N_OUT7_Mn7@263_d N_OUT6_Mn7@263_g N_VSS_Mn7@263_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@262 N_OUT7_Mn7@262_d N_OUT6_Mn7@262_g N_VSS_Mn7@262_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@263 N_OUT7_Mp7@263_d N_OUT6_Mp7@263_g N_VDD_Mp7@263_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@262 N_OUT7_Mp7@262_d N_OUT6_Mp7@262_g N_VDD_Mp7@262_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@261 N_OUT7_Mn7@261_d N_OUT6_Mn7@261_g N_VSS_Mn7@261_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@260 N_OUT7_Mn7@260_d N_OUT6_Mn7@260_g N_VSS_Mn7@260_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@261 N_OUT7_Mp7@261_d N_OUT6_Mp7@261_g N_VDD_Mp7@261_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@260 N_OUT7_Mp7@260_d N_OUT6_Mp7@260_g N_VDD_Mp7@260_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@259 N_OUT7_Mn7@259_d N_OUT6_Mn7@259_g N_VSS_Mn7@259_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@258 N_OUT7_Mn7@258_d N_OUT6_Mn7@258_g N_VSS_Mn7@258_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@259 N_OUT7_Mp7@259_d N_OUT6_Mp7@259_g N_VDD_Mp7@259_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@258 N_OUT7_Mp7@258_d N_OUT6_Mp7@258_g N_VDD_Mp7@258_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@257 N_OUT7_Mn7@257_d N_OUT6_Mn7@257_g N_VSS_Mn7@257_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@256 N_OUT7_Mn7@256_d N_OUT6_Mn7@256_g N_VSS_Mn7@256_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@257 N_OUT7_Mp7@257_d N_OUT6_Mp7@257_g N_VDD_Mp7@257_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@256 N_OUT7_Mp7@256_d N_OUT6_Mp7@256_g N_VDD_Mp7@256_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@255 N_OUT7_Mn7@255_d N_OUT6_Mn7@255_g N_VSS_Mn7@255_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@254 N_OUT7_Mn7@254_d N_OUT6_Mn7@254_g N_VSS_Mn7@254_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@255 N_OUT7_Mp7@255_d N_OUT6_Mp7@255_g N_VDD_Mp7@255_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@254 N_OUT7_Mp7@254_d N_OUT6_Mp7@254_g N_VDD_Mp7@254_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@253 N_OUT7_Mn7@253_d N_OUT6_Mn7@253_g N_VSS_Mn7@253_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@252 N_OUT7_Mn7@252_d N_OUT6_Mn7@252_g N_VSS_Mn7@252_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@253 N_OUT7_Mp7@253_d N_OUT6_Mp7@253_g N_VDD_Mp7@253_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@252 N_OUT7_Mp7@252_d N_OUT6_Mp7@252_g N_VDD_Mp7@252_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@251 N_OUT7_Mn7@251_d N_OUT6_Mn7@251_g N_VSS_Mn7@251_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@250 N_OUT7_Mn7@250_d N_OUT6_Mn7@250_g N_VSS_Mn7@250_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@251 N_OUT7_Mp7@251_d N_OUT6_Mp7@251_g N_VDD_Mp7@251_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@250 N_OUT7_Mp7@250_d N_OUT6_Mp7@250_g N_VDD_Mp7@250_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@249 N_OUT7_Mn7@249_d N_OUT6_Mn7@249_g N_VSS_Mn7@249_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@248 N_OUT7_Mn7@248_d N_OUT6_Mn7@248_g N_VSS_Mn7@248_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@249 N_OUT7_Mp7@249_d N_OUT6_Mp7@249_g N_VDD_Mp7@249_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@248 N_OUT7_Mp7@248_d N_OUT6_Mp7@248_g N_VDD_Mp7@248_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@247 N_OUT7_Mn7@247_d N_OUT6_Mn7@247_g N_VSS_Mn7@247_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@246 N_OUT7_Mn7@246_d N_OUT6_Mn7@246_g N_VSS_Mn7@246_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@247 N_OUT7_Mp7@247_d N_OUT6_Mp7@247_g N_VDD_Mp7@247_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@246 N_OUT7_Mp7@246_d N_OUT6_Mp7@246_g N_VDD_Mp7@246_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@245 N_OUT7_Mn7@245_d N_OUT6_Mn7@245_g N_VSS_Mn7@245_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@244 N_OUT7_Mn7@244_d N_OUT6_Mn7@244_g N_VSS_Mn7@244_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@245 N_OUT7_Mp7@245_d N_OUT6_Mp7@245_g N_VDD_Mp7@245_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@244 N_OUT7_Mp7@244_d N_OUT6_Mp7@244_g N_VDD_Mp7@244_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@243 N_OUT7_Mn7@243_d N_OUT6_Mn7@243_g N_VSS_Mn7@243_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@242 N_OUT7_Mn7@242_d N_OUT6_Mn7@242_g N_VSS_Mn7@242_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@243 N_OUT7_Mp7@243_d N_OUT6_Mp7@243_g N_VDD_Mp7@243_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@242 N_OUT7_Mp7@242_d N_OUT6_Mp7@242_g N_VDD_Mp7@242_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@241 N_OUT7_Mn7@241_d N_OUT6_Mn7@241_g N_VSS_Mn7@241_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@240 N_OUT7_Mn7@240_d N_OUT6_Mn7@240_g N_VSS_Mn7@240_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@241 N_OUT7_Mp7@241_d N_OUT6_Mp7@241_g N_VDD_Mp7@241_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@240 N_OUT7_Mp7@240_d N_OUT6_Mp7@240_g N_VDD_Mp7@240_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@239 N_OUT7_Mn7@239_d N_OUT6_Mn7@239_g N_VSS_Mn7@239_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@238 N_OUT7_Mn7@238_d N_OUT6_Mn7@238_g N_VSS_Mn7@238_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@239 N_OUT7_Mp7@239_d N_OUT6_Mp7@239_g N_VDD_Mp7@239_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@238 N_OUT7_Mp7@238_d N_OUT6_Mp7@238_g N_VDD_Mp7@238_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@237 N_OUT7_Mn7@237_d N_OUT6_Mn7@237_g N_VSS_Mn7@237_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@236 N_OUT7_Mn7@236_d N_OUT6_Mn7@236_g N_VSS_Mn7@236_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@237 N_OUT7_Mp7@237_d N_OUT6_Mp7@237_g N_VDD_Mp7@237_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@236 N_OUT7_Mp7@236_d N_OUT6_Mp7@236_g N_VDD_Mp7@236_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@235 N_OUT7_Mn7@235_d N_OUT6_Mn7@235_g N_VSS_Mn7@235_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@234 N_OUT7_Mn7@234_d N_OUT6_Mn7@234_g N_VSS_Mn7@234_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@235 N_OUT7_Mp7@235_d N_OUT6_Mp7@235_g N_VDD_Mp7@235_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@234 N_OUT7_Mp7@234_d N_OUT6_Mp7@234_g N_VDD_Mp7@234_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@233 N_OUT7_Mn7@233_d N_OUT6_Mn7@233_g N_VSS_Mn7@233_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@232 N_OUT7_Mn7@232_d N_OUT6_Mn7@232_g N_VSS_Mn7@232_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@233 N_OUT7_Mp7@233_d N_OUT6_Mp7@233_g N_VDD_Mp7@233_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@232 N_OUT7_Mp7@232_d N_OUT6_Mp7@232_g N_VDD_Mp7@232_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@231 N_OUT7_Mn7@231_d N_OUT6_Mn7@231_g N_VSS_Mn7@231_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@230 N_OUT7_Mn7@230_d N_OUT6_Mn7@230_g N_VSS_Mn7@230_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@231 N_OUT7_Mp7@231_d N_OUT6_Mp7@231_g N_VDD_Mp7@231_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@230 N_OUT7_Mp7@230_d N_OUT6_Mp7@230_g N_VDD_Mp7@230_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@229 N_OUT7_Mn7@229_d N_OUT6_Mn7@229_g N_VSS_Mn7@229_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@228 N_OUT7_Mn7@228_d N_OUT6_Mn7@228_g N_VSS_Mn7@228_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@229 N_OUT7_Mp7@229_d N_OUT6_Mp7@229_g N_VDD_Mp7@229_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@228 N_OUT7_Mp7@228_d N_OUT6_Mp7@228_g N_VDD_Mp7@228_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@227 N_OUT7_Mn7@227_d N_OUT6_Mn7@227_g N_VSS_Mn7@227_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@226 N_OUT7_Mn7@226_d N_OUT6_Mn7@226_g N_VSS_Mn7@226_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@227 N_OUT7_Mp7@227_d N_OUT6_Mp7@227_g N_VDD_Mp7@227_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@226 N_OUT7_Mp7@226_d N_OUT6_Mp7@226_g N_VDD_Mp7@226_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@225 N_OUT7_Mn7@225_d N_OUT6_Mn7@225_g N_VSS_Mn7@225_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@224 N_OUT7_Mn7@224_d N_OUT6_Mn7@224_g N_VSS_Mn7@224_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@225 N_OUT7_Mp7@225_d N_OUT6_Mp7@225_g N_VDD_Mp7@225_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@224 N_OUT7_Mp7@224_d N_OUT6_Mp7@224_g N_VDD_Mp7@224_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@223 N_OUT7_Mn7@223_d N_OUT6_Mn7@223_g N_VSS_Mn7@223_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@222 N_OUT7_Mn7@222_d N_OUT6_Mn7@222_g N_VSS_Mn7@222_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@223 N_OUT7_Mp7@223_d N_OUT6_Mp7@223_g N_VDD_Mp7@223_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@222 N_OUT7_Mp7@222_d N_OUT6_Mp7@222_g N_VDD_Mp7@222_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@221 N_OUT7_Mn7@221_d N_OUT6_Mn7@221_g N_VSS_Mn7@221_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@220 N_OUT7_Mn7@220_d N_OUT6_Mn7@220_g N_VSS_Mn7@220_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@221 N_OUT7_Mp7@221_d N_OUT6_Mp7@221_g N_VDD_Mp7@221_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@220 N_OUT7_Mp7@220_d N_OUT6_Mp7@220_g N_VDD_Mp7@220_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@219 N_OUT7_Mn7@219_d N_OUT6_Mn7@219_g N_VSS_Mn7@219_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@218 N_OUT7_Mn7@218_d N_OUT6_Mn7@218_g N_VSS_Mn7@218_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@219 N_OUT7_Mp7@219_d N_OUT6_Mp7@219_g N_VDD_Mp7@219_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@218 N_OUT7_Mp7@218_d N_OUT6_Mp7@218_g N_VDD_Mp7@218_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@217 N_OUT7_Mn7@217_d N_OUT6_Mn7@217_g N_VSS_Mn7@217_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@216 N_OUT7_Mn7@216_d N_OUT6_Mn7@216_g N_VSS_Mn7@216_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@217 N_OUT7_Mp7@217_d N_OUT6_Mp7@217_g N_VDD_Mp7@217_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@216 N_OUT7_Mp7@216_d N_OUT6_Mp7@216_g N_VDD_Mp7@216_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@215 N_OUT7_Mn7@215_d N_OUT6_Mn7@215_g N_VSS_Mn7@215_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@214 N_OUT7_Mn7@214_d N_OUT6_Mn7@214_g N_VSS_Mn7@214_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@215 N_OUT7_Mp7@215_d N_OUT6_Mp7@215_g N_VDD_Mp7@215_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@214 N_OUT7_Mp7@214_d N_OUT6_Mp7@214_g N_VDD_Mp7@214_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@213 N_OUT7_Mn7@213_d N_OUT6_Mn7@213_g N_VSS_Mn7@213_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@212 N_OUT7_Mn7@212_d N_OUT6_Mn7@212_g N_VSS_Mn7@212_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@213 N_OUT7_Mp7@213_d N_OUT6_Mp7@213_g N_VDD_Mp7@213_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@212 N_OUT7_Mp7@212_d N_OUT6_Mp7@212_g N_VDD_Mp7@212_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@211 N_OUT7_Mn7@211_d N_OUT6_Mn7@211_g N_VSS_Mn7@211_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@210 N_OUT7_Mn7@210_d N_OUT6_Mn7@210_g N_VSS_Mn7@210_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@211 N_OUT7_Mp7@211_d N_OUT6_Mp7@211_g N_VDD_Mp7@211_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@210 N_OUT7_Mp7@210_d N_OUT6_Mp7@210_g N_VDD_Mp7@210_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@209 N_OUT7_Mn7@209_d N_OUT6_Mn7@209_g N_VSS_Mn7@209_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@208 N_OUT7_Mn7@208_d N_OUT6_Mn7@208_g N_VSS_Mn7@208_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@209 N_OUT7_Mp7@209_d N_OUT6_Mp7@209_g N_VDD_Mp7@209_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@208 N_OUT7_Mp7@208_d N_OUT6_Mp7@208_g N_VDD_Mp7@208_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@207 N_OUT7_Mn7@207_d N_OUT6_Mn7@207_g N_VSS_Mn7@207_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@206 N_OUT7_Mn7@206_d N_OUT6_Mn7@206_g N_VSS_Mn7@206_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@207 N_OUT7_Mp7@207_d N_OUT6_Mp7@207_g N_VDD_Mp7@207_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@206 N_OUT7_Mp7@206_d N_OUT6_Mp7@206_g N_VDD_Mp7@206_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@205 N_OUT7_Mn7@205_d N_OUT6_Mn7@205_g N_VSS_Mn7@205_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@204 N_OUT7_Mn7@204_d N_OUT6_Mn7@204_g N_VSS_Mn7@204_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@205 N_OUT7_Mp7@205_d N_OUT6_Mp7@205_g N_VDD_Mp7@205_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@204 N_OUT7_Mp7@204_d N_OUT6_Mp7@204_g N_VDD_Mp7@204_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@203 N_OUT7_Mn7@203_d N_OUT6_Mn7@203_g N_VSS_Mn7@203_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@202 N_OUT7_Mn7@202_d N_OUT6_Mn7@202_g N_VSS_Mn7@202_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@203 N_OUT7_Mp7@203_d N_OUT6_Mp7@203_g N_VDD_Mp7@203_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@202 N_OUT7_Mp7@202_d N_OUT6_Mp7@202_g N_VDD_Mp7@202_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@201 N_OUT7_Mn7@201_d N_OUT6_Mn7@201_g N_VSS_Mn7@201_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@200 N_OUT7_Mn7@200_d N_OUT6_Mn7@200_g N_VSS_Mn7@200_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@201 N_OUT7_Mp7@201_d N_OUT6_Mp7@201_g N_VDD_Mp7@201_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@200 N_OUT7_Mp7@200_d N_OUT6_Mp7@200_g N_VDD_Mp7@200_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@199 N_OUT7_Mn7@199_d N_OUT6_Mn7@199_g N_VSS_Mn7@199_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@198 N_OUT7_Mn7@198_d N_OUT6_Mn7@198_g N_VSS_Mn7@198_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@199 N_OUT7_Mp7@199_d N_OUT6_Mp7@199_g N_VDD_Mp7@199_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@198 N_OUT7_Mp7@198_d N_OUT6_Mp7@198_g N_VDD_Mp7@198_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@197 N_OUT7_Mn7@197_d N_OUT6_Mn7@197_g N_VSS_Mn7@197_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@196 N_OUT7_Mn7@196_d N_OUT6_Mn7@196_g N_VSS_Mn7@196_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@197 N_OUT7_Mp7@197_d N_OUT6_Mp7@197_g N_VDD_Mp7@197_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@196 N_OUT7_Mp7@196_d N_OUT6_Mp7@196_g N_VDD_Mp7@196_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@195 N_OUT7_Mn7@195_d N_OUT6_Mn7@195_g N_VSS_Mn7@195_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@194 N_OUT7_Mn7@194_d N_OUT6_Mn7@194_g N_VSS_Mn7@194_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@195 N_OUT7_Mp7@195_d N_OUT6_Mp7@195_g N_VDD_Mp7@195_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@194 N_OUT7_Mp7@194_d N_OUT6_Mp7@194_g N_VDD_Mp7@194_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@193 N_OUT7_Mn7@193_d N_OUT6_Mn7@193_g N_VSS_Mn7@193_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@192 N_OUT7_Mn7@192_d N_OUT6_Mn7@192_g N_VSS_Mn7@192_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@193 N_OUT7_Mp7@193_d N_OUT6_Mp7@193_g N_VDD_Mp7@193_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@192 N_OUT7_Mp7@192_d N_OUT6_Mp7@192_g N_VDD_Mp7@192_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@191 N_OUT7_Mn7@191_d N_OUT6_Mn7@191_g N_VSS_Mn7@191_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@190 N_OUT7_Mn7@190_d N_OUT6_Mn7@190_g N_VSS_Mn7@190_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@191 N_OUT7_Mp7@191_d N_OUT6_Mp7@191_g N_VDD_Mp7@191_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@190 N_OUT7_Mp7@190_d N_OUT6_Mp7@190_g N_VDD_Mp7@190_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@189 N_OUT7_Mn7@189_d N_OUT6_Mn7@189_g N_VSS_Mn7@189_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@188 N_OUT7_Mn7@188_d N_OUT6_Mn7@188_g N_VSS_Mn7@188_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@189 N_OUT7_Mp7@189_d N_OUT6_Mp7@189_g N_VDD_Mp7@189_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@188 N_OUT7_Mp7@188_d N_OUT6_Mp7@188_g N_VDD_Mp7@188_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@187 N_OUT7_Mn7@187_d N_OUT6_Mn7@187_g N_VSS_Mn7@187_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@186 N_OUT7_Mn7@186_d N_OUT6_Mn7@186_g N_VSS_Mn7@186_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@187 N_OUT7_Mp7@187_d N_OUT6_Mp7@187_g N_VDD_Mp7@187_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@186 N_OUT7_Mp7@186_d N_OUT6_Mp7@186_g N_VDD_Mp7@186_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@185 N_OUT7_Mn7@185_d N_OUT6_Mn7@185_g N_VSS_Mn7@185_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@184 N_OUT7_Mn7@184_d N_OUT6_Mn7@184_g N_VSS_Mn7@184_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@185 N_OUT7_Mp7@185_d N_OUT6_Mp7@185_g N_VDD_Mp7@185_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@184 N_OUT7_Mp7@184_d N_OUT6_Mp7@184_g N_VDD_Mp7@184_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@183 N_OUT7_Mn7@183_d N_OUT6_Mn7@183_g N_VSS_Mn7@183_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@182 N_OUT7_Mn7@182_d N_OUT6_Mn7@182_g N_VSS_Mn7@182_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@183 N_OUT7_Mp7@183_d N_OUT6_Mp7@183_g N_VDD_Mp7@183_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@182 N_OUT7_Mp7@182_d N_OUT6_Mp7@182_g N_VDD_Mp7@182_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@181 N_OUT7_Mn7@181_d N_OUT6_Mn7@181_g N_VSS_Mn7@181_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@180 N_OUT7_Mn7@180_d N_OUT6_Mn7@180_g N_VSS_Mn7@180_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@181 N_OUT7_Mp7@181_d N_OUT6_Mp7@181_g N_VDD_Mp7@181_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@180 N_OUT7_Mp7@180_d N_OUT6_Mp7@180_g N_VDD_Mp7@180_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@179 N_OUT7_Mn7@179_d N_OUT6_Mn7@179_g N_VSS_Mn7@179_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@178 N_OUT7_Mn7@178_d N_OUT6_Mn7@178_g N_VSS_Mn7@178_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@179 N_OUT7_Mp7@179_d N_OUT6_Mp7@179_g N_VDD_Mp7@179_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@178 N_OUT7_Mp7@178_d N_OUT6_Mp7@178_g N_VDD_Mp7@178_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@177 N_OUT7_Mn7@177_d N_OUT6_Mn7@177_g N_VSS_Mn7@177_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@176 N_OUT7_Mn7@176_d N_OUT6_Mn7@176_g N_VSS_Mn7@176_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@177 N_OUT7_Mp7@177_d N_OUT6_Mp7@177_g N_VDD_Mp7@177_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@176 N_OUT7_Mp7@176_d N_OUT6_Mp7@176_g N_VDD_Mp7@176_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@175 N_OUT7_Mn7@175_d N_OUT6_Mn7@175_g N_VSS_Mn7@175_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@174 N_OUT7_Mn7@174_d N_OUT6_Mn7@174_g N_VSS_Mn7@174_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@175 N_OUT7_Mp7@175_d N_OUT6_Mp7@175_g N_VDD_Mp7@175_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@174 N_OUT7_Mp7@174_d N_OUT6_Mp7@174_g N_VDD_Mp7@174_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@173 N_OUT7_Mn7@173_d N_OUT6_Mn7@173_g N_VSS_Mn7@173_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@172 N_OUT7_Mn7@172_d N_OUT6_Mn7@172_g N_VSS_Mn7@172_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@173 N_OUT7_Mp7@173_d N_OUT6_Mp7@173_g N_VDD_Mp7@173_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@172 N_OUT7_Mp7@172_d N_OUT6_Mp7@172_g N_VDD_Mp7@172_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@171 N_OUT7_Mn7@171_d N_OUT6_Mn7@171_g N_VSS_Mn7@171_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@170 N_OUT7_Mn7@170_d N_OUT6_Mn7@170_g N_VSS_Mn7@170_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@171 N_OUT7_Mp7@171_d N_OUT6_Mp7@171_g N_VDD_Mp7@171_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@170 N_OUT7_Mp7@170_d N_OUT6_Mp7@170_g N_VDD_Mp7@170_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@169 N_OUT7_Mn7@169_d N_OUT6_Mn7@169_g N_VSS_Mn7@169_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@168 N_OUT7_Mn7@168_d N_OUT6_Mn7@168_g N_VSS_Mn7@168_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@169 N_OUT7_Mp7@169_d N_OUT6_Mp7@169_g N_VDD_Mp7@169_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@168 N_OUT7_Mp7@168_d N_OUT6_Mp7@168_g N_VDD_Mp7@168_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@167 N_OUT7_Mn7@167_d N_OUT6_Mn7@167_g N_VSS_Mn7@167_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@166 N_OUT7_Mn7@166_d N_OUT6_Mn7@166_g N_VSS_Mn7@166_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@167 N_OUT7_Mp7@167_d N_OUT6_Mp7@167_g N_VDD_Mp7@167_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@166 N_OUT7_Mp7@166_d N_OUT6_Mp7@166_g N_VDD_Mp7@166_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@165 N_OUT7_Mn7@165_d N_OUT6_Mn7@165_g N_VSS_Mn7@165_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@164 N_OUT7_Mn7@164_d N_OUT6_Mn7@164_g N_VSS_Mn7@164_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@165 N_OUT7_Mp7@165_d N_OUT6_Mp7@165_g N_VDD_Mp7@165_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@164 N_OUT7_Mp7@164_d N_OUT6_Mp7@164_g N_VDD_Mp7@164_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@163 N_OUT7_Mn7@163_d N_OUT6_Mn7@163_g N_VSS_Mn7@163_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@162 N_OUT7_Mn7@162_d N_OUT6_Mn7@162_g N_VSS_Mn7@162_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@163 N_OUT7_Mp7@163_d N_OUT6_Mp7@163_g N_VDD_Mp7@163_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@162 N_OUT7_Mp7@162_d N_OUT6_Mp7@162_g N_VDD_Mp7@162_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@161 N_OUT7_Mn7@161_d N_OUT6_Mn7@161_g N_VSS_Mn7@161_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@160 N_OUT7_Mn7@160_d N_OUT6_Mn7@160_g N_VSS_Mn7@160_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@161 N_OUT7_Mp7@161_d N_OUT6_Mp7@161_g N_VDD_Mp7@161_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@160 N_OUT7_Mp7@160_d N_OUT6_Mp7@160_g N_VDD_Mp7@160_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@159 N_OUT7_Mn7@159_d N_OUT6_Mn7@159_g N_VSS_Mn7@159_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@158 N_OUT7_Mn7@158_d N_OUT6_Mn7@158_g N_VSS_Mn7@158_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@159 N_OUT7_Mp7@159_d N_OUT6_Mp7@159_g N_VDD_Mp7@159_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@158 N_OUT7_Mp7@158_d N_OUT6_Mp7@158_g N_VDD_Mp7@158_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@157 N_OUT7_Mn7@157_d N_OUT6_Mn7@157_g N_VSS_Mn7@157_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@156 N_OUT7_Mn7@156_d N_OUT6_Mn7@156_g N_VSS_Mn7@156_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@157 N_OUT7_Mp7@157_d N_OUT6_Mp7@157_g N_VDD_Mp7@157_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@156 N_OUT7_Mp7@156_d N_OUT6_Mp7@156_g N_VDD_Mp7@156_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@155 N_OUT7_Mn7@155_d N_OUT6_Mn7@155_g N_VSS_Mn7@155_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@154 N_OUT7_Mn7@154_d N_OUT6_Mn7@154_g N_VSS_Mn7@154_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@155 N_OUT7_Mp7@155_d N_OUT6_Mp7@155_g N_VDD_Mp7@155_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@154 N_OUT7_Mp7@154_d N_OUT6_Mp7@154_g N_VDD_Mp7@154_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@153 N_OUT7_Mn7@153_d N_OUT6_Mn7@153_g N_VSS_Mn7@153_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@152 N_OUT7_Mn7@152_d N_OUT6_Mn7@152_g N_VSS_Mn7@152_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@153 N_OUT7_Mp7@153_d N_OUT6_Mp7@153_g N_VDD_Mp7@153_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@152 N_OUT7_Mp7@152_d N_OUT6_Mp7@152_g N_VDD_Mp7@152_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@151 N_OUT7_Mn7@151_d N_OUT6_Mn7@151_g N_VSS_Mn7@151_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@150 N_OUT7_Mn7@150_d N_OUT6_Mn7@150_g N_VSS_Mn7@150_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@151 N_OUT7_Mp7@151_d N_OUT6_Mp7@151_g N_VDD_Mp7@151_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@150 N_OUT7_Mp7@150_d N_OUT6_Mp7@150_g N_VDD_Mp7@150_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@149 N_OUT7_Mn7@149_d N_OUT6_Mn7@149_g N_VSS_Mn7@149_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@148 N_OUT7_Mn7@148_d N_OUT6_Mn7@148_g N_VSS_Mn7@148_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@149 N_OUT7_Mp7@149_d N_OUT6_Mp7@149_g N_VDD_Mp7@149_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@148 N_OUT7_Mp7@148_d N_OUT6_Mp7@148_g N_VDD_Mp7@148_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@147 N_OUT7_Mn7@147_d N_OUT6_Mn7@147_g N_VSS_Mn7@147_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@146 N_OUT7_Mn7@146_d N_OUT6_Mn7@146_g N_VSS_Mn7@146_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@147 N_OUT7_Mp7@147_d N_OUT6_Mp7@147_g N_VDD_Mp7@147_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@146 N_OUT7_Mp7@146_d N_OUT6_Mp7@146_g N_VDD_Mp7@146_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@145 N_OUT7_Mn7@145_d N_OUT6_Mn7@145_g N_VSS_Mn7@145_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@144 N_OUT7_Mn7@144_d N_OUT6_Mn7@144_g N_VSS_Mn7@144_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@145 N_OUT7_Mp7@145_d N_OUT6_Mp7@145_g N_VDD_Mp7@145_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@144 N_OUT7_Mp7@144_d N_OUT6_Mp7@144_g N_VDD_Mp7@144_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@143 N_OUT7_Mn7@143_d N_OUT6_Mn7@143_g N_VSS_Mn7@143_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@142 N_OUT7_Mn7@142_d N_OUT6_Mn7@142_g N_VSS_Mn7@142_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@143 N_OUT7_Mp7@143_d N_OUT6_Mp7@143_g N_VDD_Mp7@143_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@142 N_OUT7_Mp7@142_d N_OUT6_Mp7@142_g N_VDD_Mp7@142_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@141 N_OUT7_Mn7@141_d N_OUT6_Mn7@141_g N_VSS_Mn7@141_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@140 N_OUT7_Mn7@140_d N_OUT6_Mn7@140_g N_VSS_Mn7@140_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@141 N_OUT7_Mp7@141_d N_OUT6_Mp7@141_g N_VDD_Mp7@141_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@140 N_OUT7_Mp7@140_d N_OUT6_Mp7@140_g N_VDD_Mp7@140_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@139 N_OUT7_Mn7@139_d N_OUT6_Mn7@139_g N_VSS_Mn7@139_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@138 N_OUT7_Mn7@138_d N_OUT6_Mn7@138_g N_VSS_Mn7@138_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@139 N_OUT7_Mp7@139_d N_OUT6_Mp7@139_g N_VDD_Mp7@139_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@138 N_OUT7_Mp7@138_d N_OUT6_Mp7@138_g N_VDD_Mp7@138_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@137 N_OUT7_Mn7@137_d N_OUT6_Mn7@137_g N_VSS_Mn7@137_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@136 N_OUT7_Mn7@136_d N_OUT6_Mn7@136_g N_VSS_Mn7@136_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@137 N_OUT7_Mp7@137_d N_OUT6_Mp7@137_g N_VDD_Mp7@137_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@136 N_OUT7_Mp7@136_d N_OUT6_Mp7@136_g N_VDD_Mp7@136_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@135 N_OUT7_Mn7@135_d N_OUT6_Mn7@135_g N_VSS_Mn7@135_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@134 N_OUT7_Mn7@134_d N_OUT6_Mn7@134_g N_VSS_Mn7@134_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@135 N_OUT7_Mp7@135_d N_OUT6_Mp7@135_g N_VDD_Mp7@135_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@134 N_OUT7_Mp7@134_d N_OUT6_Mp7@134_g N_VDD_Mp7@134_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@133 N_OUT7_Mn7@133_d N_OUT6_Mn7@133_g N_VSS_Mn7@133_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@132 N_OUT7_Mn7@132_d N_OUT6_Mn7@132_g N_VSS_Mn7@132_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@133 N_OUT7_Mp7@133_d N_OUT6_Mp7@133_g N_VDD_Mp7@133_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@132 N_OUT7_Mp7@132_d N_OUT6_Mp7@132_g N_VDD_Mp7@132_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@131 N_OUT7_Mn7@131_d N_OUT6_Mn7@131_g N_VSS_Mn7@131_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@130 N_OUT7_Mn7@130_d N_OUT6_Mn7@130_g N_VSS_Mn7@130_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@131 N_OUT7_Mp7@131_d N_OUT6_Mp7@131_g N_VDD_Mp7@131_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@130 N_OUT7_Mp7@130_d N_OUT6_Mp7@130_g N_VDD_Mp7@130_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@129 N_OUT7_Mn7@129_d N_OUT6_Mn7@129_g N_VSS_Mn7@129_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@128 N_OUT7_Mn7@128_d N_OUT6_Mn7@128_g N_VSS_Mn7@128_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@129 N_OUT7_Mp7@129_d N_OUT6_Mp7@129_g N_VDD_Mp7@129_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@128 N_OUT7_Mp7@128_d N_OUT6_Mp7@128_g N_VDD_Mp7@128_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@127 N_OUT7_Mn7@127_d N_OUT6_Mn7@127_g N_VSS_Mn7@127_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@126 N_OUT7_Mn7@126_d N_OUT6_Mn7@126_g N_VSS_Mn7@126_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@127 N_OUT7_Mp7@127_d N_OUT6_Mp7@127_g N_VDD_Mp7@127_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@126 N_OUT7_Mp7@126_d N_OUT6_Mp7@126_g N_VDD_Mp7@126_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@125 N_OUT7_Mn7@125_d N_OUT6_Mn7@125_g N_VSS_Mn7@125_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@124 N_OUT7_Mn7@124_d N_OUT6_Mn7@124_g N_VSS_Mn7@124_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@125 N_OUT7_Mp7@125_d N_OUT6_Mp7@125_g N_VDD_Mp7@125_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@124 N_OUT7_Mp7@124_d N_OUT6_Mp7@124_g N_VDD_Mp7@124_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@123 N_OUT7_Mn7@123_d N_OUT6_Mn7@123_g N_VSS_Mn7@123_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@122 N_OUT7_Mn7@122_d N_OUT6_Mn7@122_g N_VSS_Mn7@122_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@123 N_OUT7_Mp7@123_d N_OUT6_Mp7@123_g N_VDD_Mp7@123_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@122 N_OUT7_Mp7@122_d N_OUT6_Mp7@122_g N_VDD_Mp7@122_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@121 N_OUT7_Mn7@121_d N_OUT6_Mn7@121_g N_VSS_Mn7@121_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@120 N_OUT7_Mn7@120_d N_OUT6_Mn7@120_g N_VSS_Mn7@120_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@121 N_OUT7_Mp7@121_d N_OUT6_Mp7@121_g N_VDD_Mp7@121_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@120 N_OUT7_Mp7@120_d N_OUT6_Mp7@120_g N_VDD_Mp7@120_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@119 N_OUT7_Mn7@119_d N_OUT6_Mn7@119_g N_VSS_Mn7@119_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@118 N_OUT7_Mn7@118_d N_OUT6_Mn7@118_g N_VSS_Mn7@118_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@119 N_OUT7_Mp7@119_d N_OUT6_Mp7@119_g N_VDD_Mp7@119_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@118 N_OUT7_Mp7@118_d N_OUT6_Mp7@118_g N_VDD_Mp7@118_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@117 N_OUT7_Mn7@117_d N_OUT6_Mn7@117_g N_VSS_Mn7@117_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@116 N_OUT7_Mn7@116_d N_OUT6_Mn7@116_g N_VSS_Mn7@116_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@117 N_OUT7_Mp7@117_d N_OUT6_Mp7@117_g N_VDD_Mp7@117_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@116 N_OUT7_Mp7@116_d N_OUT6_Mp7@116_g N_VDD_Mp7@116_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@115 N_OUT7_Mn7@115_d N_OUT6_Mn7@115_g N_VSS_Mn7@115_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@114 N_OUT7_Mn7@114_d N_OUT6_Mn7@114_g N_VSS_Mn7@114_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@115 N_OUT7_Mp7@115_d N_OUT6_Mp7@115_g N_VDD_Mp7@115_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@114 N_OUT7_Mp7@114_d N_OUT6_Mp7@114_g N_VDD_Mp7@114_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@113 N_OUT7_Mn7@113_d N_OUT6_Mn7@113_g N_VSS_Mn7@113_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@112 N_OUT7_Mn7@112_d N_OUT6_Mn7@112_g N_VSS_Mn7@112_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@113 N_OUT7_Mp7@113_d N_OUT6_Mp7@113_g N_VDD_Mp7@113_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@112 N_OUT7_Mp7@112_d N_OUT6_Mp7@112_g N_VDD_Mp7@112_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@111 N_OUT7_Mn7@111_d N_OUT6_Mn7@111_g N_VSS_Mn7@111_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@110 N_OUT7_Mn7@110_d N_OUT6_Mn7@110_g N_VSS_Mn7@110_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@111 N_OUT7_Mp7@111_d N_OUT6_Mp7@111_g N_VDD_Mp7@111_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@110 N_OUT7_Mp7@110_d N_OUT6_Mp7@110_g N_VDD_Mp7@110_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@109 N_OUT7_Mn7@109_d N_OUT6_Mn7@109_g N_VSS_Mn7@109_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@108 N_OUT7_Mn7@108_d N_OUT6_Mn7@108_g N_VSS_Mn7@108_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@109 N_OUT7_Mp7@109_d N_OUT6_Mp7@109_g N_VDD_Mp7@109_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@108 N_OUT7_Mp7@108_d N_OUT6_Mp7@108_g N_VDD_Mp7@108_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@107 N_OUT7_Mn7@107_d N_OUT6_Mn7@107_g N_VSS_Mn7@107_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@106 N_OUT7_Mn7@106_d N_OUT6_Mn7@106_g N_VSS_Mn7@106_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@107 N_OUT7_Mp7@107_d N_OUT6_Mp7@107_g N_VDD_Mp7@107_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@106 N_OUT7_Mp7@106_d N_OUT6_Mp7@106_g N_VDD_Mp7@106_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@105 N_OUT7_Mn7@105_d N_OUT6_Mn7@105_g N_VSS_Mn7@105_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@104 N_OUT7_Mn7@104_d N_OUT6_Mn7@104_g N_VSS_Mn7@104_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@105 N_OUT7_Mp7@105_d N_OUT6_Mp7@105_g N_VDD_Mp7@105_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@104 N_OUT7_Mp7@104_d N_OUT6_Mp7@104_g N_VDD_Mp7@104_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@103 N_OUT7_Mn7@103_d N_OUT6_Mn7@103_g N_VSS_Mn7@103_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@102 N_OUT7_Mn7@102_d N_OUT6_Mn7@102_g N_VSS_Mn7@102_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@103 N_OUT7_Mp7@103_d N_OUT6_Mp7@103_g N_VDD_Mp7@103_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@102 N_OUT7_Mp7@102_d N_OUT6_Mp7@102_g N_VDD_Mp7@102_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@101 N_OUT7_Mn7@101_d N_OUT6_Mn7@101_g N_VSS_Mn7@101_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@100 N_OUT7_Mn7@100_d N_OUT6_Mn7@100_g N_VSS_Mn7@100_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@101 N_OUT7_Mp7@101_d N_OUT6_Mp7@101_g N_VDD_Mp7@101_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@100 N_OUT7_Mp7@100_d N_OUT6_Mp7@100_g N_VDD_Mp7@100_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@99 N_OUT7_Mn7@99_d N_OUT6_Mn7@99_g N_VSS_Mn7@99_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@98 N_OUT7_Mn7@98_d N_OUT6_Mn7@98_g N_VSS_Mn7@98_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@99 N_OUT7_Mp7@99_d N_OUT6_Mp7@99_g N_VDD_Mp7@99_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@98 N_OUT7_Mp7@98_d N_OUT6_Mp7@98_g N_VDD_Mp7@98_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@97 N_OUT7_Mn7@97_d N_OUT6_Mn7@97_g N_VSS_Mn7@97_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@96 N_OUT7_Mn7@96_d N_OUT6_Mn7@96_g N_VSS_Mn7@96_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@97 N_OUT7_Mp7@97_d N_OUT6_Mp7@97_g N_VDD_Mp7@97_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@96 N_OUT7_Mp7@96_d N_OUT6_Mp7@96_g N_VDD_Mp7@96_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@95 N_OUT7_Mn7@95_d N_OUT6_Mn7@95_g N_VSS_Mn7@95_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@94 N_OUT7_Mn7@94_d N_OUT6_Mn7@94_g N_VSS_Mn7@94_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@95 N_OUT7_Mp7@95_d N_OUT6_Mp7@95_g N_VDD_Mp7@95_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@94 N_OUT7_Mp7@94_d N_OUT6_Mp7@94_g N_VDD_Mp7@94_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@93 N_OUT7_Mn7@93_d N_OUT6_Mn7@93_g N_VSS_Mn7@93_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@92 N_OUT7_Mn7@92_d N_OUT6_Mn7@92_g N_VSS_Mn7@92_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@93 N_OUT7_Mp7@93_d N_OUT6_Mp7@93_g N_VDD_Mp7@93_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@92 N_OUT7_Mp7@92_d N_OUT6_Mp7@92_g N_VDD_Mp7@92_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@91 N_OUT7_Mn7@91_d N_OUT6_Mn7@91_g N_VSS_Mn7@91_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@90 N_OUT7_Mn7@90_d N_OUT6_Mn7@90_g N_VSS_Mn7@90_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@91 N_OUT7_Mp7@91_d N_OUT6_Mp7@91_g N_VDD_Mp7@91_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@90 N_OUT7_Mp7@90_d N_OUT6_Mp7@90_g N_VDD_Mp7@90_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@89 N_OUT7_Mn7@89_d N_OUT6_Mn7@89_g N_VSS_Mn7@89_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@88 N_OUT7_Mn7@88_d N_OUT6_Mn7@88_g N_VSS_Mn7@88_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@89 N_OUT7_Mp7@89_d N_OUT6_Mp7@89_g N_VDD_Mp7@89_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@88 N_OUT7_Mp7@88_d N_OUT6_Mp7@88_g N_VDD_Mp7@88_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@87 N_OUT7_Mn7@87_d N_OUT6_Mn7@87_g N_VSS_Mn7@87_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@86 N_OUT7_Mn7@86_d N_OUT6_Mn7@86_g N_VSS_Mn7@86_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@87 N_OUT7_Mp7@87_d N_OUT6_Mp7@87_g N_VDD_Mp7@87_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@86 N_OUT7_Mp7@86_d N_OUT6_Mp7@86_g N_VDD_Mp7@86_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@85 N_OUT7_Mn7@85_d N_OUT6_Mn7@85_g N_VSS_Mn7@85_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@84 N_OUT7_Mn7@84_d N_OUT6_Mn7@84_g N_VSS_Mn7@84_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@85 N_OUT7_Mp7@85_d N_OUT6_Mp7@85_g N_VDD_Mp7@85_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@84 N_OUT7_Mp7@84_d N_OUT6_Mp7@84_g N_VDD_Mp7@84_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@83 N_OUT7_Mn7@83_d N_OUT6_Mn7@83_g N_VSS_Mn7@83_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@82 N_OUT7_Mn7@82_d N_OUT6_Mn7@82_g N_VSS_Mn7@82_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@83 N_OUT7_Mp7@83_d N_OUT6_Mp7@83_g N_VDD_Mp7@83_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@82 N_OUT7_Mp7@82_d N_OUT6_Mp7@82_g N_VDD_Mp7@82_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@81 N_OUT7_Mn7@81_d N_OUT6_Mn7@81_g N_VSS_Mn7@81_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@80 N_OUT7_Mn7@80_d N_OUT6_Mn7@80_g N_VSS_Mn7@80_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@81 N_OUT7_Mp7@81_d N_OUT6_Mp7@81_g N_VDD_Mp7@81_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@80 N_OUT7_Mp7@80_d N_OUT6_Mp7@80_g N_VDD_Mp7@80_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@79 N_OUT7_Mn7@79_d N_OUT6_Mn7@79_g N_VSS_Mn7@79_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@78 N_OUT7_Mn7@78_d N_OUT6_Mn7@78_g N_VSS_Mn7@78_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@79 N_OUT7_Mp7@79_d N_OUT6_Mp7@79_g N_VDD_Mp7@79_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@78 N_OUT7_Mp7@78_d N_OUT6_Mp7@78_g N_VDD_Mp7@78_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@77 N_OUT7_Mn7@77_d N_OUT6_Mn7@77_g N_VSS_Mn7@77_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@76 N_OUT7_Mn7@76_d N_OUT6_Mn7@76_g N_VSS_Mn7@76_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@77 N_OUT7_Mp7@77_d N_OUT6_Mp7@77_g N_VDD_Mp7@77_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@76 N_OUT7_Mp7@76_d N_OUT6_Mp7@76_g N_VDD_Mp7@76_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@75 N_OUT7_Mn7@75_d N_OUT6_Mn7@75_g N_VSS_Mn7@75_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@74 N_OUT7_Mn7@74_d N_OUT6_Mn7@74_g N_VSS_Mn7@74_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@75 N_OUT7_Mp7@75_d N_OUT6_Mp7@75_g N_VDD_Mp7@75_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@74 N_OUT7_Mp7@74_d N_OUT6_Mp7@74_g N_VDD_Mp7@74_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@73 N_OUT7_Mn7@73_d N_OUT6_Mn7@73_g N_VSS_Mn7@73_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@72 N_OUT7_Mn7@72_d N_OUT6_Mn7@72_g N_VSS_Mn7@72_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@73 N_OUT7_Mp7@73_d N_OUT6_Mp7@73_g N_VDD_Mp7@73_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@72 N_OUT7_Mp7@72_d N_OUT6_Mp7@72_g N_VDD_Mp7@72_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@71 N_OUT7_Mn7@71_d N_OUT6_Mn7@71_g N_VSS_Mn7@71_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@70 N_OUT7_Mn7@70_d N_OUT6_Mn7@70_g N_VSS_Mn7@70_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@71 N_OUT7_Mp7@71_d N_OUT6_Mp7@71_g N_VDD_Mp7@71_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@70 N_OUT7_Mp7@70_d N_OUT6_Mp7@70_g N_VDD_Mp7@70_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@69 N_OUT7_Mn7@69_d N_OUT6_Mn7@69_g N_VSS_Mn7@69_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@68 N_OUT7_Mn7@68_d N_OUT6_Mn7@68_g N_VSS_Mn7@68_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@69 N_OUT7_Mp7@69_d N_OUT6_Mp7@69_g N_VDD_Mp7@69_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@68 N_OUT7_Mp7@68_d N_OUT6_Mp7@68_g N_VDD_Mp7@68_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@67 N_OUT7_Mn7@67_d N_OUT6_Mn7@67_g N_VSS_Mn7@67_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@66 N_OUT7_Mn7@66_d N_OUT6_Mn7@66_g N_VSS_Mn7@66_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@67 N_OUT7_Mp7@67_d N_OUT6_Mp7@67_g N_VDD_Mp7@67_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@66 N_OUT7_Mp7@66_d N_OUT6_Mp7@66_g N_VDD_Mp7@66_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@65 N_OUT7_Mn7@65_d N_OUT6_Mn7@65_g N_VSS_Mn7@65_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@64 N_OUT7_Mn7@64_d N_OUT6_Mn7@64_g N_VSS_Mn7@64_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@65 N_OUT7_Mp7@65_d N_OUT6_Mp7@65_g N_VDD_Mp7@65_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@64 N_OUT7_Mp7@64_d N_OUT6_Mp7@64_g N_VDD_Mp7@64_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@63 N_OUT7_Mn7@63_d N_OUT6_Mn7@63_g N_VSS_Mn7@63_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@62 N_OUT7_Mn7@62_d N_OUT6_Mn7@62_g N_VSS_Mn7@62_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@63 N_OUT7_Mp7@63_d N_OUT6_Mp7@63_g N_VDD_Mp7@63_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@62 N_OUT7_Mp7@62_d N_OUT6_Mp7@62_g N_VDD_Mp7@62_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@61 N_OUT7_Mn7@61_d N_OUT6_Mn7@61_g N_VSS_Mn7@61_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@60 N_OUT7_Mn7@60_d N_OUT6_Mn7@60_g N_VSS_Mn7@60_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@61 N_OUT7_Mp7@61_d N_OUT6_Mp7@61_g N_VDD_Mp7@61_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@60 N_OUT7_Mp7@60_d N_OUT6_Mp7@60_g N_VDD_Mp7@60_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@59 N_OUT7_Mn7@59_d N_OUT6_Mn7@59_g N_VSS_Mn7@59_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@58 N_OUT7_Mn7@58_d N_OUT6_Mn7@58_g N_VSS_Mn7@58_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@59 N_OUT7_Mp7@59_d N_OUT6_Mp7@59_g N_VDD_Mp7@59_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@58 N_OUT7_Mp7@58_d N_OUT6_Mp7@58_g N_VDD_Mp7@58_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@57 N_OUT7_Mn7@57_d N_OUT6_Mn7@57_g N_VSS_Mn7@57_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@56 N_OUT7_Mn7@56_d N_OUT6_Mn7@56_g N_VSS_Mn7@56_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@57 N_OUT7_Mp7@57_d N_OUT6_Mp7@57_g N_VDD_Mp7@57_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@56 N_OUT7_Mp7@56_d N_OUT6_Mp7@56_g N_VDD_Mp7@56_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@55 N_OUT7_Mn7@55_d N_OUT6_Mn7@55_g N_VSS_Mn7@55_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@54 N_OUT7_Mn7@54_d N_OUT6_Mn7@54_g N_VSS_Mn7@54_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@55 N_OUT7_Mp7@55_d N_OUT6_Mp7@55_g N_VDD_Mp7@55_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@54 N_OUT7_Mp7@54_d N_OUT6_Mp7@54_g N_VDD_Mp7@54_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@53 N_OUT7_Mn7@53_d N_OUT6_Mn7@53_g N_VSS_Mn7@53_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@52 N_OUT7_Mn7@52_d N_OUT6_Mn7@52_g N_VSS_Mn7@52_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@53 N_OUT7_Mp7@53_d N_OUT6_Mp7@53_g N_VDD_Mp7@53_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@52 N_OUT7_Mp7@52_d N_OUT6_Mp7@52_g N_VDD_Mp7@52_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@51 N_OUT7_Mn7@51_d N_OUT6_Mn7@51_g N_VSS_Mn7@51_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@50 N_OUT7_Mn7@50_d N_OUT6_Mn7@50_g N_VSS_Mn7@50_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@51 N_OUT7_Mp7@51_d N_OUT6_Mp7@51_g N_VDD_Mp7@51_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@50 N_OUT7_Mp7@50_d N_OUT6_Mp7@50_g N_VDD_Mp7@50_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@49 N_OUT7_Mn7@49_d N_OUT6_Mn7@49_g N_VSS_Mn7@49_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@48 N_OUT7_Mn7@48_d N_OUT6_Mn7@48_g N_VSS_Mn7@48_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@49 N_OUT7_Mp7@49_d N_OUT6_Mp7@49_g N_VDD_Mp7@49_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@48 N_OUT7_Mp7@48_d N_OUT6_Mp7@48_g N_VDD_Mp7@48_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@47 N_OUT7_Mn7@47_d N_OUT6_Mn7@47_g N_VSS_Mn7@47_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@46 N_OUT7_Mn7@46_d N_OUT6_Mn7@46_g N_VSS_Mn7@46_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@47 N_OUT7_Mp7@47_d N_OUT6_Mp7@47_g N_VDD_Mp7@47_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@46 N_OUT7_Mp7@46_d N_OUT6_Mp7@46_g N_VDD_Mp7@46_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@45 N_OUT7_Mn7@45_d N_OUT6_Mn7@45_g N_VSS_Mn7@45_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@44 N_OUT7_Mn7@44_d N_OUT6_Mn7@44_g N_VSS_Mn7@44_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@45 N_OUT7_Mp7@45_d N_OUT6_Mp7@45_g N_VDD_Mp7@45_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@44 N_OUT7_Mp7@44_d N_OUT6_Mp7@44_g N_VDD_Mp7@44_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@43 N_OUT7_Mn7@43_d N_OUT6_Mn7@43_g N_VSS_Mn7@43_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@42 N_OUT7_Mn7@42_d N_OUT6_Mn7@42_g N_VSS_Mn7@42_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@43 N_OUT7_Mp7@43_d N_OUT6_Mp7@43_g N_VDD_Mp7@43_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@42 N_OUT7_Mp7@42_d N_OUT6_Mp7@42_g N_VDD_Mp7@42_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@41 N_OUT7_Mn7@41_d N_OUT6_Mn7@41_g N_VSS_Mn7@41_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@40 N_OUT7_Mn7@40_d N_OUT6_Mn7@40_g N_VSS_Mn7@40_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@41 N_OUT7_Mp7@41_d N_OUT6_Mp7@41_g N_VDD_Mp7@41_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@40 N_OUT7_Mp7@40_d N_OUT6_Mp7@40_g N_VDD_Mp7@40_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@39 N_OUT7_Mn7@39_d N_OUT6_Mn7@39_g N_VSS_Mn7@39_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@38 N_OUT7_Mn7@38_d N_OUT6_Mn7@38_g N_VSS_Mn7@38_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@39 N_OUT7_Mp7@39_d N_OUT6_Mp7@39_g N_VDD_Mp7@39_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@38 N_OUT7_Mp7@38_d N_OUT6_Mp7@38_g N_VDD_Mp7@38_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@37 N_OUT7_Mn7@37_d N_OUT6_Mn7@37_g N_VSS_Mn7@37_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@36 N_OUT7_Mn7@36_d N_OUT6_Mn7@36_g N_VSS_Mn7@36_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@37 N_OUT7_Mp7@37_d N_OUT6_Mp7@37_g N_VDD_Mp7@37_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@36 N_OUT7_Mp7@36_d N_OUT6_Mp7@36_g N_VDD_Mp7@36_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@35 N_OUT7_Mn7@35_d N_OUT6_Mn7@35_g N_VSS_Mn7@35_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@34 N_OUT7_Mn7@34_d N_OUT6_Mn7@34_g N_VSS_Mn7@34_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@35 N_OUT7_Mp7@35_d N_OUT6_Mp7@35_g N_VDD_Mp7@35_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@34 N_OUT7_Mp7@34_d N_OUT6_Mp7@34_g N_VDD_Mp7@34_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@33 N_OUT7_Mn7@33_d N_OUT6_Mn7@33_g N_VSS_Mn7@33_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@32 N_OUT7_Mn7@32_d N_OUT6_Mn7@32_g N_VSS_Mn7@32_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@33 N_OUT7_Mp7@33_d N_OUT6_Mp7@33_g N_VDD_Mp7@33_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@32 N_OUT7_Mp7@32_d N_OUT6_Mp7@32_g N_VDD_Mp7@32_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@31 N_OUT7_Mn7@31_d N_OUT6_Mn7@31_g N_VSS_Mn7@31_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@30 N_OUT7_Mn7@30_d N_OUT6_Mn7@30_g N_VSS_Mn7@30_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@31 N_OUT7_Mp7@31_d N_OUT6_Mp7@31_g N_VDD_Mp7@31_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@30 N_OUT7_Mp7@30_d N_OUT6_Mp7@30_g N_VDD_Mp7@30_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@29 N_OUT7_Mn7@29_d N_OUT6_Mn7@29_g N_VSS_Mn7@29_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@28 N_OUT7_Mn7@28_d N_OUT6_Mn7@28_g N_VSS_Mn7@28_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@29 N_OUT7_Mp7@29_d N_OUT6_Mp7@29_g N_VDD_Mp7@29_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@28 N_OUT7_Mp7@28_d N_OUT6_Mp7@28_g N_VDD_Mp7@28_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@27 N_OUT7_Mn7@27_d N_OUT6_Mn7@27_g N_VSS_Mn7@27_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@26 N_OUT7_Mn7@26_d N_OUT6_Mn7@26_g N_VSS_Mn7@26_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@27 N_OUT7_Mp7@27_d N_OUT6_Mp7@27_g N_VDD_Mp7@27_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@26 N_OUT7_Mp7@26_d N_OUT6_Mp7@26_g N_VDD_Mp7@26_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@25 N_OUT7_Mn7@25_d N_OUT6_Mn7@25_g N_VSS_Mn7@25_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@24 N_OUT7_Mn7@24_d N_OUT6_Mn7@24_g N_VSS_Mn7@24_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@25 N_OUT7_Mp7@25_d N_OUT6_Mp7@25_g N_VDD_Mp7@25_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@24 N_OUT7_Mp7@24_d N_OUT6_Mp7@24_g N_VDD_Mp7@24_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@23 N_OUT7_Mn7@23_d N_OUT6_Mn7@23_g N_VSS_Mn7@23_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@22 N_OUT7_Mn7@22_d N_OUT6_Mn7@22_g N_VSS_Mn7@22_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@23 N_OUT7_Mp7@23_d N_OUT6_Mp7@23_g N_VDD_Mp7@23_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@22 N_OUT7_Mp7@22_d N_OUT6_Mp7@22_g N_VDD_Mp7@22_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@21 N_OUT7_Mn7@21_d N_OUT6_Mn7@21_g N_VSS_Mn7@21_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@20 N_OUT7_Mn7@20_d N_OUT6_Mn7@20_g N_VSS_Mn7@20_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@21 N_OUT7_Mp7@21_d N_OUT6_Mp7@21_g N_VDD_Mp7@21_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@20 N_OUT7_Mp7@20_d N_OUT6_Mp7@20_g N_VDD_Mp7@20_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@19 N_OUT7_Mn7@19_d N_OUT6_Mn7@19_g N_VSS_Mn7@19_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@18 N_OUT7_Mn7@18_d N_OUT6_Mn7@18_g N_VSS_Mn7@18_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@19 N_OUT7_Mp7@19_d N_OUT6_Mp7@19_g N_VDD_Mp7@19_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@18 N_OUT7_Mp7@18_d N_OUT6_Mp7@18_g N_VDD_Mp7@18_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@17 N_OUT7_Mn7@17_d N_OUT6_Mn7@17_g N_VSS_Mn7@17_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@16 N_OUT7_Mn7@16_d N_OUT6_Mn7@16_g N_VSS_Mn7@16_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@17 N_OUT7_Mp7@17_d N_OUT6_Mp7@17_g N_VDD_Mp7@17_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@16 N_OUT7_Mp7@16_d N_OUT6_Mp7@16_g N_VDD_Mp7@16_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@15 N_OUT7_Mn7@15_d N_OUT6_Mn7@15_g N_VSS_Mn7@15_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@14 N_OUT7_Mn7@14_d N_OUT6_Mn7@14_g N_VSS_Mn7@14_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@15 N_OUT7_Mp7@15_d N_OUT6_Mp7@15_g N_VDD_Mp7@15_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@14 N_OUT7_Mp7@14_d N_OUT6_Mp7@14_g N_VDD_Mp7@14_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@13 N_OUT7_Mn7@13_d N_OUT6_Mn7@13_g N_VSS_Mn7@13_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@12 N_OUT7_Mn7@12_d N_OUT6_Mn7@12_g N_VSS_Mn7@12_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@13 N_OUT7_Mp7@13_d N_OUT6_Mp7@13_g N_VDD_Mp7@13_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@12 N_OUT7_Mp7@12_d N_OUT6_Mp7@12_g N_VDD_Mp7@12_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@11 N_OUT7_Mn7@11_d N_OUT6_Mn7@11_g N_VSS_Mn7@11_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@10 N_OUT7_Mn7@10_d N_OUT6_Mn7@10_g N_VSS_Mn7@10_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@11 N_OUT7_Mp7@11_d N_OUT6_Mp7@11_g N_VDD_Mp7@11_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@10 N_OUT7_Mp7@10_d N_OUT6_Mp7@10_g N_VDD_Mp7@10_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@9 N_OUT7_Mn7@9_d N_OUT6_Mn7@9_g N_VSS_Mn7@9_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@8 N_OUT7_Mn7@8_d N_OUT6_Mn7@8_g N_VSS_Mn7@8_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@9 N_OUT7_Mp7@9_d N_OUT6_Mp7@9_g N_VDD_Mp7@9_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@8 N_OUT7_Mp7@8_d N_OUT6_Mp7@8_g N_VDD_Mp7@8_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@7 N_OUT7_Mn7@7_d N_OUT6_Mn7@7_g N_VSS_Mn7@7_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@6 N_OUT7_Mn7@6_d N_OUT6_Mn7@6_g N_VSS_Mn7@6_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@7 N_OUT7_Mp7@7_d N_OUT6_Mp7@7_g N_VDD_Mp7@7_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@6 N_OUT7_Mp7@6_d N_OUT6_Mp7@6_g N_VDD_Mp7@6_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@5 N_OUT7_Mn7@5_d N_OUT6_Mn7@5_g N_VSS_Mn7@5_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@4 N_OUT7_Mn7@4_d N_OUT6_Mn7@4_g N_VSS_Mn7@4_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@5 N_OUT7_Mp7@5_d N_OUT6_Mp7@5_g N_VDD_Mp7@5_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@4 N_OUT7_Mp7@4_d N_OUT6_Mp7@4_g N_VDD_Mp7@4_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn7@3 N_OUT7_Mn7@3_d N_OUT6_Mn7@3_g N_VSS_Mn7@3_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn7@2 N_OUT7_Mn7@2_d N_OUT6_Mn7@2_g N_VSS_Mn7@2_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp7@3 N_OUT7_Mp7@3_d N_OUT6_Mp7@3_g N_VDD_Mp7@3_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp7@2 N_OUT7_Mp7@2_d N_OUT6_Mp7@2_g N_VDD_Mp7@2_s N_VDD_Mp7@1159_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3073 N_OUT8_Mn8@3073_d N_OUT7_Mn8@3073_g N_VSS_Mn8@3073_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3072 N_OUT8_Mn8@3072_d N_OUT7_Mn8@3072_g N_VSS_Mn8@3072_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3073 N_OUT8_Mp8@3073_d N_OUT7_Mp8@3073_g N_VDD_Mp8@3073_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3072 N_OUT8_Mp8@3072_d N_OUT7_Mp8@3072_g N_VDD_Mp8@3072_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3071 N_OUT8_Mn8@3071_d N_OUT7_Mn8@3071_g N_VSS_Mn8@3071_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3070 N_OUT8_Mn8@3070_d N_OUT7_Mn8@3070_g N_VSS_Mn8@3070_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3071 N_OUT8_Mp8@3071_d N_OUT7_Mp8@3071_g N_VDD_Mp8@3071_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3070 N_OUT8_Mp8@3070_d N_OUT7_Mp8@3070_g N_VDD_Mp8@3070_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3069 N_OUT8_Mn8@3069_d N_OUT7_Mn8@3069_g N_VSS_Mn8@3069_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3068 N_OUT8_Mn8@3068_d N_OUT7_Mn8@3068_g N_VSS_Mn8@3068_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3069 N_OUT8_Mp8@3069_d N_OUT7_Mp8@3069_g N_VDD_Mp8@3069_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3068 N_OUT8_Mp8@3068_d N_OUT7_Mp8@3068_g N_VDD_Mp8@3068_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3067 N_OUT8_Mn8@3067_d N_OUT7_Mn8@3067_g N_VSS_Mn8@3067_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3066 N_OUT8_Mn8@3066_d N_OUT7_Mn8@3066_g N_VSS_Mn8@3066_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3067 N_OUT8_Mp8@3067_d N_OUT7_Mp8@3067_g N_VDD_Mp8@3067_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3066 N_OUT8_Mp8@3066_d N_OUT7_Mp8@3066_g N_VDD_Mp8@3066_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3065 N_OUT8_Mn8@3065_d N_OUT7_Mn8@3065_g N_VSS_Mn8@3065_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3064 N_OUT8_Mn8@3064_d N_OUT7_Mn8@3064_g N_VSS_Mn8@3064_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3065 N_OUT8_Mp8@3065_d N_OUT7_Mp8@3065_g N_VDD_Mp8@3065_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3064 N_OUT8_Mp8@3064_d N_OUT7_Mp8@3064_g N_VDD_Mp8@3064_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3063 N_OUT8_Mn8@3063_d N_OUT7_Mn8@3063_g N_VSS_Mn8@3063_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3062 N_OUT8_Mn8@3062_d N_OUT7_Mn8@3062_g N_VSS_Mn8@3062_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3063 N_OUT8_Mp8@3063_d N_OUT7_Mp8@3063_g N_VDD_Mp8@3063_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3062 N_OUT8_Mp8@3062_d N_OUT7_Mp8@3062_g N_VDD_Mp8@3062_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3061 N_OUT8_Mn8@3061_d N_OUT7_Mn8@3061_g N_VSS_Mn8@3061_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3060 N_OUT8_Mn8@3060_d N_OUT7_Mn8@3060_g N_VSS_Mn8@3060_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3061 N_OUT8_Mp8@3061_d N_OUT7_Mp8@3061_g N_VDD_Mp8@3061_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3060 N_OUT8_Mp8@3060_d N_OUT7_Mp8@3060_g N_VDD_Mp8@3060_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3059 N_OUT8_Mn8@3059_d N_OUT7_Mn8@3059_g N_VSS_Mn8@3059_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3058 N_OUT8_Mn8@3058_d N_OUT7_Mn8@3058_g N_VSS_Mn8@3058_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3059 N_OUT8_Mp8@3059_d N_OUT7_Mp8@3059_g N_VDD_Mp8@3059_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3058 N_OUT8_Mp8@3058_d N_OUT7_Mp8@3058_g N_VDD_Mp8@3058_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3057 N_OUT8_Mn8@3057_d N_OUT7_Mn8@3057_g N_VSS_Mn8@3057_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3056 N_OUT8_Mn8@3056_d N_OUT7_Mn8@3056_g N_VSS_Mn8@3056_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3057 N_OUT8_Mp8@3057_d N_OUT7_Mp8@3057_g N_VDD_Mp8@3057_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3056 N_OUT8_Mp8@3056_d N_OUT7_Mp8@3056_g N_VDD_Mp8@3056_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3055 N_OUT8_Mn8@3055_d N_OUT7_Mn8@3055_g N_VSS_Mn8@3055_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3054 N_OUT8_Mn8@3054_d N_OUT7_Mn8@3054_g N_VSS_Mn8@3054_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3055 N_OUT8_Mp8@3055_d N_OUT7_Mp8@3055_g N_VDD_Mp8@3055_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3054 N_OUT8_Mp8@3054_d N_OUT7_Mp8@3054_g N_VDD_Mp8@3054_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3053 N_OUT8_Mn8@3053_d N_OUT7_Mn8@3053_g N_VSS_Mn8@3053_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3052 N_OUT8_Mn8@3052_d N_OUT7_Mn8@3052_g N_VSS_Mn8@3052_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3053 N_OUT8_Mp8@3053_d N_OUT7_Mp8@3053_g N_VDD_Mp8@3053_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3052 N_OUT8_Mp8@3052_d N_OUT7_Mp8@3052_g N_VDD_Mp8@3052_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3051 N_OUT8_Mn8@3051_d N_OUT7_Mn8@3051_g N_VSS_Mn8@3051_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3050 N_OUT8_Mn8@3050_d N_OUT7_Mn8@3050_g N_VSS_Mn8@3050_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3051 N_OUT8_Mp8@3051_d N_OUT7_Mp8@3051_g N_VDD_Mp8@3051_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3050 N_OUT8_Mp8@3050_d N_OUT7_Mp8@3050_g N_VDD_Mp8@3050_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3049 N_OUT8_Mn8@3049_d N_OUT7_Mn8@3049_g N_VSS_Mn8@3049_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3048 N_OUT8_Mn8@3048_d N_OUT7_Mn8@3048_g N_VSS_Mn8@3048_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3049 N_OUT8_Mp8@3049_d N_OUT7_Mp8@3049_g N_VDD_Mp8@3049_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3048 N_OUT8_Mp8@3048_d N_OUT7_Mp8@3048_g N_VDD_Mp8@3048_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3047 N_OUT8_Mn8@3047_d N_OUT7_Mn8@3047_g N_VSS_Mn8@3047_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3046 N_OUT8_Mn8@3046_d N_OUT7_Mn8@3046_g N_VSS_Mn8@3046_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3047 N_OUT8_Mp8@3047_d N_OUT7_Mp8@3047_g N_VDD_Mp8@3047_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3046 N_OUT8_Mp8@3046_d N_OUT7_Mp8@3046_g N_VDD_Mp8@3046_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3045 N_OUT8_Mn8@3045_d N_OUT7_Mn8@3045_g N_VSS_Mn8@3045_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3044 N_OUT8_Mn8@3044_d N_OUT7_Mn8@3044_g N_VSS_Mn8@3044_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3045 N_OUT8_Mp8@3045_d N_OUT7_Mp8@3045_g N_VDD_Mp8@3045_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3044 N_OUT8_Mp8@3044_d N_OUT7_Mp8@3044_g N_VDD_Mp8@3044_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3043 N_OUT8_Mn8@3043_d N_OUT7_Mn8@3043_g N_VSS_Mn8@3043_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3042 N_OUT8_Mn8@3042_d N_OUT7_Mn8@3042_g N_VSS_Mn8@3042_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3043 N_OUT8_Mp8@3043_d N_OUT7_Mp8@3043_g N_VDD_Mp8@3043_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3042 N_OUT8_Mp8@3042_d N_OUT7_Mp8@3042_g N_VDD_Mp8@3042_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3041 N_OUT8_Mn8@3041_d N_OUT7_Mn8@3041_g N_VSS_Mn8@3041_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3040 N_OUT8_Mn8@3040_d N_OUT7_Mn8@3040_g N_VSS_Mn8@3040_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3041 N_OUT8_Mp8@3041_d N_OUT7_Mp8@3041_g N_VDD_Mp8@3041_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3040 N_OUT8_Mp8@3040_d N_OUT7_Mp8@3040_g N_VDD_Mp8@3040_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3039 N_OUT8_Mn8@3039_d N_OUT7_Mn8@3039_g N_VSS_Mn8@3039_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3038 N_OUT8_Mn8@3038_d N_OUT7_Mn8@3038_g N_VSS_Mn8@3038_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3039 N_OUT8_Mp8@3039_d N_OUT7_Mp8@3039_g N_VDD_Mp8@3039_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3038 N_OUT8_Mp8@3038_d N_OUT7_Mp8@3038_g N_VDD_Mp8@3038_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3037 N_OUT8_Mn8@3037_d N_OUT7_Mn8@3037_g N_VSS_Mn8@3037_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3036 N_OUT8_Mn8@3036_d N_OUT7_Mn8@3036_g N_VSS_Mn8@3036_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3037 N_OUT8_Mp8@3037_d N_OUT7_Mp8@3037_g N_VDD_Mp8@3037_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3036 N_OUT8_Mp8@3036_d N_OUT7_Mp8@3036_g N_VDD_Mp8@3036_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3035 N_OUT8_Mn8@3035_d N_OUT7_Mn8@3035_g N_VSS_Mn8@3035_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3034 N_OUT8_Mn8@3034_d N_OUT7_Mn8@3034_g N_VSS_Mn8@3034_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3035 N_OUT8_Mp8@3035_d N_OUT7_Mp8@3035_g N_VDD_Mp8@3035_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3034 N_OUT8_Mp8@3034_d N_OUT7_Mp8@3034_g N_VDD_Mp8@3034_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3033 N_OUT8_Mn8@3033_d N_OUT7_Mn8@3033_g N_VSS_Mn8@3033_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3032 N_OUT8_Mn8@3032_d N_OUT7_Mn8@3032_g N_VSS_Mn8@3032_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3033 N_OUT8_Mp8@3033_d N_OUT7_Mp8@3033_g N_VDD_Mp8@3033_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3032 N_OUT8_Mp8@3032_d N_OUT7_Mp8@3032_g N_VDD_Mp8@3032_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3031 N_OUT8_Mn8@3031_d N_OUT7_Mn8@3031_g N_VSS_Mn8@3031_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3030 N_OUT8_Mn8@3030_d N_OUT7_Mn8@3030_g N_VSS_Mn8@3030_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3031 N_OUT8_Mp8@3031_d N_OUT7_Mp8@3031_g N_VDD_Mp8@3031_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3030 N_OUT8_Mp8@3030_d N_OUT7_Mp8@3030_g N_VDD_Mp8@3030_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3029 N_OUT8_Mn8@3029_d N_OUT7_Mn8@3029_g N_VSS_Mn8@3029_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3028 N_OUT8_Mn8@3028_d N_OUT7_Mn8@3028_g N_VSS_Mn8@3028_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3029 N_OUT8_Mp8@3029_d N_OUT7_Mp8@3029_g N_VDD_Mp8@3029_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3028 N_OUT8_Mp8@3028_d N_OUT7_Mp8@3028_g N_VDD_Mp8@3028_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3027 N_OUT8_Mn8@3027_d N_OUT7_Mn8@3027_g N_VSS_Mn8@3027_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3026 N_OUT8_Mn8@3026_d N_OUT7_Mn8@3026_g N_VSS_Mn8@3026_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3027 N_OUT8_Mp8@3027_d N_OUT7_Mp8@3027_g N_VDD_Mp8@3027_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3026 N_OUT8_Mp8@3026_d N_OUT7_Mp8@3026_g N_VDD_Mp8@3026_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3025 N_OUT8_Mn8@3025_d N_OUT7_Mn8@3025_g N_VSS_Mn8@3025_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3024 N_OUT8_Mn8@3024_d N_OUT7_Mn8@3024_g N_VSS_Mn8@3024_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3025 N_OUT8_Mp8@3025_d N_OUT7_Mp8@3025_g N_VDD_Mp8@3025_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3024 N_OUT8_Mp8@3024_d N_OUT7_Mp8@3024_g N_VDD_Mp8@3024_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3023 N_OUT8_Mn8@3023_d N_OUT7_Mn8@3023_g N_VSS_Mn8@3023_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3022 N_OUT8_Mn8@3022_d N_OUT7_Mn8@3022_g N_VSS_Mn8@3022_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3023 N_OUT8_Mp8@3023_d N_OUT7_Mp8@3023_g N_VDD_Mp8@3023_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3022 N_OUT8_Mp8@3022_d N_OUT7_Mp8@3022_g N_VDD_Mp8@3022_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3021 N_OUT8_Mn8@3021_d N_OUT7_Mn8@3021_g N_VSS_Mn8@3021_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3020 N_OUT8_Mn8@3020_d N_OUT7_Mn8@3020_g N_VSS_Mn8@3020_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3021 N_OUT8_Mp8@3021_d N_OUT7_Mp8@3021_g N_VDD_Mp8@3021_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3020 N_OUT8_Mp8@3020_d N_OUT7_Mp8@3020_g N_VDD_Mp8@3020_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3019 N_OUT8_Mn8@3019_d N_OUT7_Mn8@3019_g N_VSS_Mn8@3019_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3018 N_OUT8_Mn8@3018_d N_OUT7_Mn8@3018_g N_VSS_Mn8@3018_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3019 N_OUT8_Mp8@3019_d N_OUT7_Mp8@3019_g N_VDD_Mp8@3019_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3018 N_OUT8_Mp8@3018_d N_OUT7_Mp8@3018_g N_VDD_Mp8@3018_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3017 N_OUT8_Mn8@3017_d N_OUT7_Mn8@3017_g N_VSS_Mn8@3017_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3016 N_OUT8_Mn8@3016_d N_OUT7_Mn8@3016_g N_VSS_Mn8@3016_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3017 N_OUT8_Mp8@3017_d N_OUT7_Mp8@3017_g N_VDD_Mp8@3017_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3016 N_OUT8_Mp8@3016_d N_OUT7_Mp8@3016_g N_VDD_Mp8@3016_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3015 N_OUT8_Mn8@3015_d N_OUT7_Mn8@3015_g N_VSS_Mn8@3015_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3014 N_OUT8_Mn8@3014_d N_OUT7_Mn8@3014_g N_VSS_Mn8@3014_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3015 N_OUT8_Mp8@3015_d N_OUT7_Mp8@3015_g N_VDD_Mp8@3015_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3014 N_OUT8_Mp8@3014_d N_OUT7_Mp8@3014_g N_VDD_Mp8@3014_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3013 N_OUT8_Mn8@3013_d N_OUT7_Mn8@3013_g N_VSS_Mn8@3013_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3012 N_OUT8_Mn8@3012_d N_OUT7_Mn8@3012_g N_VSS_Mn8@3012_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3013 N_OUT8_Mp8@3013_d N_OUT7_Mp8@3013_g N_VDD_Mp8@3013_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3012 N_OUT8_Mp8@3012_d N_OUT7_Mp8@3012_g N_VDD_Mp8@3012_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3011 N_OUT8_Mn8@3011_d N_OUT7_Mn8@3011_g N_VSS_Mn8@3011_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3010 N_OUT8_Mn8@3010_d N_OUT7_Mn8@3010_g N_VSS_Mn8@3010_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3011 N_OUT8_Mp8@3011_d N_OUT7_Mp8@3011_g N_VDD_Mp8@3011_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3010 N_OUT8_Mp8@3010_d N_OUT7_Mp8@3010_g N_VDD_Mp8@3010_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3009 N_OUT8_Mn8@3009_d N_OUT7_Mn8@3009_g N_VSS_Mn8@3009_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3008 N_OUT8_Mn8@3008_d N_OUT7_Mn8@3008_g N_VSS_Mn8@3008_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3009 N_OUT8_Mp8@3009_d N_OUT7_Mp8@3009_g N_VDD_Mp8@3009_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3008 N_OUT8_Mp8@3008_d N_OUT7_Mp8@3008_g N_VDD_Mp8@3008_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3007 N_OUT8_Mn8@3007_d N_OUT7_Mn8@3007_g N_VSS_Mn8@3007_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3006 N_OUT8_Mn8@3006_d N_OUT7_Mn8@3006_g N_VSS_Mn8@3006_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3007 N_OUT8_Mp8@3007_d N_OUT7_Mp8@3007_g N_VDD_Mp8@3007_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3006 N_OUT8_Mp8@3006_d N_OUT7_Mp8@3006_g N_VDD_Mp8@3006_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3005 N_OUT8_Mn8@3005_d N_OUT7_Mn8@3005_g N_VSS_Mn8@3005_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3004 N_OUT8_Mn8@3004_d N_OUT7_Mn8@3004_g N_VSS_Mn8@3004_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3005 N_OUT8_Mp8@3005_d N_OUT7_Mp8@3005_g N_VDD_Mp8@3005_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3004 N_OUT8_Mp8@3004_d N_OUT7_Mp8@3004_g N_VDD_Mp8@3004_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3003 N_OUT8_Mn8@3003_d N_OUT7_Mn8@3003_g N_VSS_Mn8@3003_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3002 N_OUT8_Mn8@3002_d N_OUT7_Mn8@3002_g N_VSS_Mn8@3002_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3003 N_OUT8_Mp8@3003_d N_OUT7_Mp8@3003_g N_VDD_Mp8@3003_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3002 N_OUT8_Mp8@3002_d N_OUT7_Mp8@3002_g N_VDD_Mp8@3002_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3001 N_OUT8_Mn8@3001_d N_OUT7_Mn8@3001_g N_VSS_Mn8@3001_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@3000 N_OUT8_Mn8@3000_d N_OUT7_Mn8@3000_g N_VSS_Mn8@3000_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3001 N_OUT8_Mp8@3001_d N_OUT7_Mp8@3001_g N_VDD_Mp8@3001_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@3000 N_OUT8_Mp8@3000_d N_OUT7_Mp8@3000_g N_VDD_Mp8@3000_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2999 N_OUT8_Mn8@2999_d N_OUT7_Mn8@2999_g N_VSS_Mn8@2999_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2998 N_OUT8_Mn8@2998_d N_OUT7_Mn8@2998_g N_VSS_Mn8@2998_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2999 N_OUT8_Mp8@2999_d N_OUT7_Mp8@2999_g N_VDD_Mp8@2999_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2998 N_OUT8_Mp8@2998_d N_OUT7_Mp8@2998_g N_VDD_Mp8@2998_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2997 N_OUT8_Mn8@2997_d N_OUT7_Mn8@2997_g N_VSS_Mn8@2997_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2996 N_OUT8_Mn8@2996_d N_OUT7_Mn8@2996_g N_VSS_Mn8@2996_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2997 N_OUT8_Mp8@2997_d N_OUT7_Mp8@2997_g N_VDD_Mp8@2997_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2996 N_OUT8_Mp8@2996_d N_OUT7_Mp8@2996_g N_VDD_Mp8@2996_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2995 N_OUT8_Mn8@2995_d N_OUT7_Mn8@2995_g N_VSS_Mn8@2995_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2994 N_OUT8_Mn8@2994_d N_OUT7_Mn8@2994_g N_VSS_Mn8@2994_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2995 N_OUT8_Mp8@2995_d N_OUT7_Mp8@2995_g N_VDD_Mp8@2995_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2994 N_OUT8_Mp8@2994_d N_OUT7_Mp8@2994_g N_VDD_Mp8@2994_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2993 N_OUT8_Mn8@2993_d N_OUT7_Mn8@2993_g N_VSS_Mn8@2993_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2992 N_OUT8_Mn8@2992_d N_OUT7_Mn8@2992_g N_VSS_Mn8@2992_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2993 N_OUT8_Mp8@2993_d N_OUT7_Mp8@2993_g N_VDD_Mp8@2993_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2992 N_OUT8_Mp8@2992_d N_OUT7_Mp8@2992_g N_VDD_Mp8@2992_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2991 N_OUT8_Mn8@2991_d N_OUT7_Mn8@2991_g N_VSS_Mn8@2991_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2990 N_OUT8_Mn8@2990_d N_OUT7_Mn8@2990_g N_VSS_Mn8@2990_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2991 N_OUT8_Mp8@2991_d N_OUT7_Mp8@2991_g N_VDD_Mp8@2991_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2990 N_OUT8_Mp8@2990_d N_OUT7_Mp8@2990_g N_VDD_Mp8@2990_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2989 N_OUT8_Mn8@2989_d N_OUT7_Mn8@2989_g N_VSS_Mn8@2989_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2988 N_OUT8_Mn8@2988_d N_OUT7_Mn8@2988_g N_VSS_Mn8@2988_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2989 N_OUT8_Mp8@2989_d N_OUT7_Mp8@2989_g N_VDD_Mp8@2989_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2988 N_OUT8_Mp8@2988_d N_OUT7_Mp8@2988_g N_VDD_Mp8@2988_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2987 N_OUT8_Mn8@2987_d N_OUT7_Mn8@2987_g N_VSS_Mn8@2987_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2986 N_OUT8_Mn8@2986_d N_OUT7_Mn8@2986_g N_VSS_Mn8@2986_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2987 N_OUT8_Mp8@2987_d N_OUT7_Mp8@2987_g N_VDD_Mp8@2987_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2986 N_OUT8_Mp8@2986_d N_OUT7_Mp8@2986_g N_VDD_Mp8@2986_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2985 N_OUT8_Mn8@2985_d N_OUT7_Mn8@2985_g N_VSS_Mn8@2985_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2984 N_OUT8_Mn8@2984_d N_OUT7_Mn8@2984_g N_VSS_Mn8@2984_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2985 N_OUT8_Mp8@2985_d N_OUT7_Mp8@2985_g N_VDD_Mp8@2985_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2984 N_OUT8_Mp8@2984_d N_OUT7_Mp8@2984_g N_VDD_Mp8@2984_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2983 N_OUT8_Mn8@2983_d N_OUT7_Mn8@2983_g N_VSS_Mn8@2983_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2982 N_OUT8_Mn8@2982_d N_OUT7_Mn8@2982_g N_VSS_Mn8@2982_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2983 N_OUT8_Mp8@2983_d N_OUT7_Mp8@2983_g N_VDD_Mp8@2983_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2982 N_OUT8_Mp8@2982_d N_OUT7_Mp8@2982_g N_VDD_Mp8@2982_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2981 N_OUT8_Mn8@2981_d N_OUT7_Mn8@2981_g N_VSS_Mn8@2981_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2980 N_OUT8_Mn8@2980_d N_OUT7_Mn8@2980_g N_VSS_Mn8@2980_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2981 N_OUT8_Mp8@2981_d N_OUT7_Mp8@2981_g N_VDD_Mp8@2981_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2980 N_OUT8_Mp8@2980_d N_OUT7_Mp8@2980_g N_VDD_Mp8@2980_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2979 N_OUT8_Mn8@2979_d N_OUT7_Mn8@2979_g N_VSS_Mn8@2979_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2978 N_OUT8_Mn8@2978_d N_OUT7_Mn8@2978_g N_VSS_Mn8@2978_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2979 N_OUT8_Mp8@2979_d N_OUT7_Mp8@2979_g N_VDD_Mp8@2979_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2978 N_OUT8_Mp8@2978_d N_OUT7_Mp8@2978_g N_VDD_Mp8@2978_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2977 N_OUT8_Mn8@2977_d N_OUT7_Mn8@2977_g N_VSS_Mn8@2977_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2976 N_OUT8_Mn8@2976_d N_OUT7_Mn8@2976_g N_VSS_Mn8@2976_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2977 N_OUT8_Mp8@2977_d N_OUT7_Mp8@2977_g N_VDD_Mp8@2977_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2976 N_OUT8_Mp8@2976_d N_OUT7_Mp8@2976_g N_VDD_Mp8@2976_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2975 N_OUT8_Mn8@2975_d N_OUT7_Mn8@2975_g N_VSS_Mn8@2975_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2974 N_OUT8_Mn8@2974_d N_OUT7_Mn8@2974_g N_VSS_Mn8@2974_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2975 N_OUT8_Mp8@2975_d N_OUT7_Mp8@2975_g N_VDD_Mp8@2975_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2974 N_OUT8_Mp8@2974_d N_OUT7_Mp8@2974_g N_VDD_Mp8@2974_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2973 N_OUT8_Mn8@2973_d N_OUT7_Mn8@2973_g N_VSS_Mn8@2973_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2972 N_OUT8_Mn8@2972_d N_OUT7_Mn8@2972_g N_VSS_Mn8@2972_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2973 N_OUT8_Mp8@2973_d N_OUT7_Mp8@2973_g N_VDD_Mp8@2973_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2972 N_OUT8_Mp8@2972_d N_OUT7_Mp8@2972_g N_VDD_Mp8@2972_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2971 N_OUT8_Mn8@2971_d N_OUT7_Mn8@2971_g N_VSS_Mn8@2971_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2970 N_OUT8_Mn8@2970_d N_OUT7_Mn8@2970_g N_VSS_Mn8@2970_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2971 N_OUT8_Mp8@2971_d N_OUT7_Mp8@2971_g N_VDD_Mp8@2971_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2970 N_OUT8_Mp8@2970_d N_OUT7_Mp8@2970_g N_VDD_Mp8@2970_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2969 N_OUT8_Mn8@2969_d N_OUT7_Mn8@2969_g N_VSS_Mn8@2969_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2968 N_OUT8_Mn8@2968_d N_OUT7_Mn8@2968_g N_VSS_Mn8@2968_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2969 N_OUT8_Mp8@2969_d N_OUT7_Mp8@2969_g N_VDD_Mp8@2969_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2968 N_OUT8_Mp8@2968_d N_OUT7_Mp8@2968_g N_VDD_Mp8@2968_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2967 N_OUT8_Mn8@2967_d N_OUT7_Mn8@2967_g N_VSS_Mn8@2967_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2966 N_OUT8_Mn8@2966_d N_OUT7_Mn8@2966_g N_VSS_Mn8@2966_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2967 N_OUT8_Mp8@2967_d N_OUT7_Mp8@2967_g N_VDD_Mp8@2967_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2966 N_OUT8_Mp8@2966_d N_OUT7_Mp8@2966_g N_VDD_Mp8@2966_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2965 N_OUT8_Mn8@2965_d N_OUT7_Mn8@2965_g N_VSS_Mn8@2965_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2964 N_OUT8_Mn8@2964_d N_OUT7_Mn8@2964_g N_VSS_Mn8@2964_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2965 N_OUT8_Mp8@2965_d N_OUT7_Mp8@2965_g N_VDD_Mp8@2965_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2964 N_OUT8_Mp8@2964_d N_OUT7_Mp8@2964_g N_VDD_Mp8@2964_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2963 N_OUT8_Mn8@2963_d N_OUT7_Mn8@2963_g N_VSS_Mn8@2963_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2962 N_OUT8_Mn8@2962_d N_OUT7_Mn8@2962_g N_VSS_Mn8@2962_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2963 N_OUT8_Mp8@2963_d N_OUT7_Mp8@2963_g N_VDD_Mp8@2963_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2962 N_OUT8_Mp8@2962_d N_OUT7_Mp8@2962_g N_VDD_Mp8@2962_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2961 N_OUT8_Mn8@2961_d N_OUT7_Mn8@2961_g N_VSS_Mn8@2961_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2960 N_OUT8_Mn8@2960_d N_OUT7_Mn8@2960_g N_VSS_Mn8@2960_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2961 N_OUT8_Mp8@2961_d N_OUT7_Mp8@2961_g N_VDD_Mp8@2961_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2960 N_OUT8_Mp8@2960_d N_OUT7_Mp8@2960_g N_VDD_Mp8@2960_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2959 N_OUT8_Mn8@2959_d N_OUT7_Mn8@2959_g N_VSS_Mn8@2959_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2958 N_OUT8_Mn8@2958_d N_OUT7_Mn8@2958_g N_VSS_Mn8@2958_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2959 N_OUT8_Mp8@2959_d N_OUT7_Mp8@2959_g N_VDD_Mp8@2959_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2958 N_OUT8_Mp8@2958_d N_OUT7_Mp8@2958_g N_VDD_Mp8@2958_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2957 N_OUT8_Mn8@2957_d N_OUT7_Mn8@2957_g N_VSS_Mn8@2957_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2956 N_OUT8_Mn8@2956_d N_OUT7_Mn8@2956_g N_VSS_Mn8@2956_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2957 N_OUT8_Mp8@2957_d N_OUT7_Mp8@2957_g N_VDD_Mp8@2957_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2956 N_OUT8_Mp8@2956_d N_OUT7_Mp8@2956_g N_VDD_Mp8@2956_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2955 N_OUT8_Mn8@2955_d N_OUT7_Mn8@2955_g N_VSS_Mn8@2955_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2954 N_OUT8_Mn8@2954_d N_OUT7_Mn8@2954_g N_VSS_Mn8@2954_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2955 N_OUT8_Mp8@2955_d N_OUT7_Mp8@2955_g N_VDD_Mp8@2955_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2954 N_OUT8_Mp8@2954_d N_OUT7_Mp8@2954_g N_VDD_Mp8@2954_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2953 N_OUT8_Mn8@2953_d N_OUT7_Mn8@2953_g N_VSS_Mn8@2953_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2952 N_OUT8_Mn8@2952_d N_OUT7_Mn8@2952_g N_VSS_Mn8@2952_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2953 N_OUT8_Mp8@2953_d N_OUT7_Mp8@2953_g N_VDD_Mp8@2953_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2952 N_OUT8_Mp8@2952_d N_OUT7_Mp8@2952_g N_VDD_Mp8@2952_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2951 N_OUT8_Mn8@2951_d N_OUT7_Mn8@2951_g N_VSS_Mn8@2951_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2950 N_OUT8_Mn8@2950_d N_OUT7_Mn8@2950_g N_VSS_Mn8@2950_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2951 N_OUT8_Mp8@2951_d N_OUT7_Mp8@2951_g N_VDD_Mp8@2951_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2950 N_OUT8_Mp8@2950_d N_OUT7_Mp8@2950_g N_VDD_Mp8@2950_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2949 N_OUT8_Mn8@2949_d N_OUT7_Mn8@2949_g N_VSS_Mn8@2949_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2948 N_OUT8_Mn8@2948_d N_OUT7_Mn8@2948_g N_VSS_Mn8@2948_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2949 N_OUT8_Mp8@2949_d N_OUT7_Mp8@2949_g N_VDD_Mp8@2949_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2948 N_OUT8_Mp8@2948_d N_OUT7_Mp8@2948_g N_VDD_Mp8@2948_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2947 N_OUT8_Mn8@2947_d N_OUT7_Mn8@2947_g N_VSS_Mn8@2947_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2946 N_OUT8_Mn8@2946_d N_OUT7_Mn8@2946_g N_VSS_Mn8@2946_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2947 N_OUT8_Mp8@2947_d N_OUT7_Mp8@2947_g N_VDD_Mp8@2947_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2946 N_OUT8_Mp8@2946_d N_OUT7_Mp8@2946_g N_VDD_Mp8@2946_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2945 N_OUT8_Mn8@2945_d N_OUT7_Mn8@2945_g N_VSS_Mn8@2945_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2944 N_OUT8_Mn8@2944_d N_OUT7_Mn8@2944_g N_VSS_Mn8@2944_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2945 N_OUT8_Mp8@2945_d N_OUT7_Mp8@2945_g N_VDD_Mp8@2945_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2944 N_OUT8_Mp8@2944_d N_OUT7_Mp8@2944_g N_VDD_Mp8@2944_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2943 N_OUT8_Mn8@2943_d N_OUT7_Mn8@2943_g N_VSS_Mn8@2943_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2942 N_OUT8_Mn8@2942_d N_OUT7_Mn8@2942_g N_VSS_Mn8@2942_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2943 N_OUT8_Mp8@2943_d N_OUT7_Mp8@2943_g N_VDD_Mp8@2943_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2942 N_OUT8_Mp8@2942_d N_OUT7_Mp8@2942_g N_VDD_Mp8@2942_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2941 N_OUT8_Mn8@2941_d N_OUT7_Mn8@2941_g N_VSS_Mn8@2941_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2940 N_OUT8_Mn8@2940_d N_OUT7_Mn8@2940_g N_VSS_Mn8@2940_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2941 N_OUT8_Mp8@2941_d N_OUT7_Mp8@2941_g N_VDD_Mp8@2941_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2940 N_OUT8_Mp8@2940_d N_OUT7_Mp8@2940_g N_VDD_Mp8@2940_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2939 N_OUT8_Mn8@2939_d N_OUT7_Mn8@2939_g N_VSS_Mn8@2939_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2938 N_OUT8_Mn8@2938_d N_OUT7_Mn8@2938_g N_VSS_Mn8@2938_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2939 N_OUT8_Mp8@2939_d N_OUT7_Mp8@2939_g N_VDD_Mp8@2939_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2938 N_OUT8_Mp8@2938_d N_OUT7_Mp8@2938_g N_VDD_Mp8@2938_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2937 N_OUT8_Mn8@2937_d N_OUT7_Mn8@2937_g N_VSS_Mn8@2937_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2936 N_OUT8_Mn8@2936_d N_OUT7_Mn8@2936_g N_VSS_Mn8@2936_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2937 N_OUT8_Mp8@2937_d N_OUT7_Mp8@2937_g N_VDD_Mp8@2937_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2936 N_OUT8_Mp8@2936_d N_OUT7_Mp8@2936_g N_VDD_Mp8@2936_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2935 N_OUT8_Mn8@2935_d N_OUT7_Mn8@2935_g N_VSS_Mn8@2935_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2934 N_OUT8_Mn8@2934_d N_OUT7_Mn8@2934_g N_VSS_Mn8@2934_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2935 N_OUT8_Mp8@2935_d N_OUT7_Mp8@2935_g N_VDD_Mp8@2935_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2934 N_OUT8_Mp8@2934_d N_OUT7_Mp8@2934_g N_VDD_Mp8@2934_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2933 N_OUT8_Mn8@2933_d N_OUT7_Mn8@2933_g N_VSS_Mn8@2933_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2932 N_OUT8_Mn8@2932_d N_OUT7_Mn8@2932_g N_VSS_Mn8@2932_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2933 N_OUT8_Mp8@2933_d N_OUT7_Mp8@2933_g N_VDD_Mp8@2933_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2932 N_OUT8_Mp8@2932_d N_OUT7_Mp8@2932_g N_VDD_Mp8@2932_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2931 N_OUT8_Mn8@2931_d N_OUT7_Mn8@2931_g N_VSS_Mn8@2931_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2930 N_OUT8_Mn8@2930_d N_OUT7_Mn8@2930_g N_VSS_Mn8@2930_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2931 N_OUT8_Mp8@2931_d N_OUT7_Mp8@2931_g N_VDD_Mp8@2931_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2930 N_OUT8_Mp8@2930_d N_OUT7_Mp8@2930_g N_VDD_Mp8@2930_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2929 N_OUT8_Mn8@2929_d N_OUT7_Mn8@2929_g N_VSS_Mn8@2929_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2928 N_OUT8_Mn8@2928_d N_OUT7_Mn8@2928_g N_VSS_Mn8@2928_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2929 N_OUT8_Mp8@2929_d N_OUT7_Mp8@2929_g N_VDD_Mp8@2929_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2928 N_OUT8_Mp8@2928_d N_OUT7_Mp8@2928_g N_VDD_Mp8@2928_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2927 N_OUT8_Mn8@2927_d N_OUT7_Mn8@2927_g N_VSS_Mn8@2927_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2926 N_OUT8_Mn8@2926_d N_OUT7_Mn8@2926_g N_VSS_Mn8@2926_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2927 N_OUT8_Mp8@2927_d N_OUT7_Mp8@2927_g N_VDD_Mp8@2927_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2926 N_OUT8_Mp8@2926_d N_OUT7_Mp8@2926_g N_VDD_Mp8@2926_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2925 N_OUT8_Mn8@2925_d N_OUT7_Mn8@2925_g N_VSS_Mn8@2925_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2924 N_OUT8_Mn8@2924_d N_OUT7_Mn8@2924_g N_VSS_Mn8@2924_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2925 N_OUT8_Mp8@2925_d N_OUT7_Mp8@2925_g N_VDD_Mp8@2925_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2924 N_OUT8_Mp8@2924_d N_OUT7_Mp8@2924_g N_VDD_Mp8@2924_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2923 N_OUT8_Mn8@2923_d N_OUT7_Mn8@2923_g N_VSS_Mn8@2923_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2922 N_OUT8_Mn8@2922_d N_OUT7_Mn8@2922_g N_VSS_Mn8@2922_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2923 N_OUT8_Mp8@2923_d N_OUT7_Mp8@2923_g N_VDD_Mp8@2923_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2922 N_OUT8_Mp8@2922_d N_OUT7_Mp8@2922_g N_VDD_Mp8@2922_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2921 N_OUT8_Mn8@2921_d N_OUT7_Mn8@2921_g N_VSS_Mn8@2921_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2920 N_OUT8_Mn8@2920_d N_OUT7_Mn8@2920_g N_VSS_Mn8@2920_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2921 N_OUT8_Mp8@2921_d N_OUT7_Mp8@2921_g N_VDD_Mp8@2921_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2920 N_OUT8_Mp8@2920_d N_OUT7_Mp8@2920_g N_VDD_Mp8@2920_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2919 N_OUT8_Mn8@2919_d N_OUT7_Mn8@2919_g N_VSS_Mn8@2919_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2918 N_OUT8_Mn8@2918_d N_OUT7_Mn8@2918_g N_VSS_Mn8@2918_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2919 N_OUT8_Mp8@2919_d N_OUT7_Mp8@2919_g N_VDD_Mp8@2919_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2918 N_OUT8_Mp8@2918_d N_OUT7_Mp8@2918_g N_VDD_Mp8@2918_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2917 N_OUT8_Mn8@2917_d N_OUT7_Mn8@2917_g N_VSS_Mn8@2917_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2916 N_OUT8_Mn8@2916_d N_OUT7_Mn8@2916_g N_VSS_Mn8@2916_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2917 N_OUT8_Mp8@2917_d N_OUT7_Mp8@2917_g N_VDD_Mp8@2917_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2916 N_OUT8_Mp8@2916_d N_OUT7_Mp8@2916_g N_VDD_Mp8@2916_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2915 N_OUT8_Mn8@2915_d N_OUT7_Mn8@2915_g N_VSS_Mn8@2915_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2914 N_OUT8_Mn8@2914_d N_OUT7_Mn8@2914_g N_VSS_Mn8@2914_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2915 N_OUT8_Mp8@2915_d N_OUT7_Mp8@2915_g N_VDD_Mp8@2915_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2914 N_OUT8_Mp8@2914_d N_OUT7_Mp8@2914_g N_VDD_Mp8@2914_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2913 N_OUT8_Mn8@2913_d N_OUT7_Mn8@2913_g N_VSS_Mn8@2913_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2912 N_OUT8_Mn8@2912_d N_OUT7_Mn8@2912_g N_VSS_Mn8@2912_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2913 N_OUT8_Mp8@2913_d N_OUT7_Mp8@2913_g N_VDD_Mp8@2913_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2912 N_OUT8_Mp8@2912_d N_OUT7_Mp8@2912_g N_VDD_Mp8@2912_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2911 N_OUT8_Mn8@2911_d N_OUT7_Mn8@2911_g N_VSS_Mn8@2911_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2910 N_OUT8_Mn8@2910_d N_OUT7_Mn8@2910_g N_VSS_Mn8@2910_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2911 N_OUT8_Mp8@2911_d N_OUT7_Mp8@2911_g N_VDD_Mp8@2911_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2910 N_OUT8_Mp8@2910_d N_OUT7_Mp8@2910_g N_VDD_Mp8@2910_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2909 N_OUT8_Mn8@2909_d N_OUT7_Mn8@2909_g N_VSS_Mn8@2909_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2908 N_OUT8_Mn8@2908_d N_OUT7_Mn8@2908_g N_VSS_Mn8@2908_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2909 N_OUT8_Mp8@2909_d N_OUT7_Mp8@2909_g N_VDD_Mp8@2909_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2908 N_OUT8_Mp8@2908_d N_OUT7_Mp8@2908_g N_VDD_Mp8@2908_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2907 N_OUT8_Mn8@2907_d N_OUT7_Mn8@2907_g N_VSS_Mn8@2907_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2906 N_OUT8_Mn8@2906_d N_OUT7_Mn8@2906_g N_VSS_Mn8@2906_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2907 N_OUT8_Mp8@2907_d N_OUT7_Mp8@2907_g N_VDD_Mp8@2907_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2906 N_OUT8_Mp8@2906_d N_OUT7_Mp8@2906_g N_VDD_Mp8@2906_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2905 N_OUT8_Mn8@2905_d N_OUT7_Mn8@2905_g N_VSS_Mn8@2905_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2904 N_OUT8_Mn8@2904_d N_OUT7_Mn8@2904_g N_VSS_Mn8@2904_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2905 N_OUT8_Mp8@2905_d N_OUT7_Mp8@2905_g N_VDD_Mp8@2905_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2904 N_OUT8_Mp8@2904_d N_OUT7_Mp8@2904_g N_VDD_Mp8@2904_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2903 N_OUT8_Mn8@2903_d N_OUT7_Mn8@2903_g N_VSS_Mn8@2903_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2902 N_OUT8_Mn8@2902_d N_OUT7_Mn8@2902_g N_VSS_Mn8@2902_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2903 N_OUT8_Mp8@2903_d N_OUT7_Mp8@2903_g N_VDD_Mp8@2903_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2902 N_OUT8_Mp8@2902_d N_OUT7_Mp8@2902_g N_VDD_Mp8@2902_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2901 N_OUT8_Mn8@2901_d N_OUT7_Mn8@2901_g N_VSS_Mn8@2901_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2900 N_OUT8_Mn8@2900_d N_OUT7_Mn8@2900_g N_VSS_Mn8@2900_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2901 N_OUT8_Mp8@2901_d N_OUT7_Mp8@2901_g N_VDD_Mp8@2901_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2900 N_OUT8_Mp8@2900_d N_OUT7_Mp8@2900_g N_VDD_Mp8@2900_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2899 N_OUT8_Mn8@2899_d N_OUT7_Mn8@2899_g N_VSS_Mn8@2899_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2898 N_OUT8_Mn8@2898_d N_OUT7_Mn8@2898_g N_VSS_Mn8@2898_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2899 N_OUT8_Mp8@2899_d N_OUT7_Mp8@2899_g N_VDD_Mp8@2899_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2898 N_OUT8_Mp8@2898_d N_OUT7_Mp8@2898_g N_VDD_Mp8@2898_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2897 N_OUT8_Mn8@2897_d N_OUT7_Mn8@2897_g N_VSS_Mn8@2897_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2896 N_OUT8_Mn8@2896_d N_OUT7_Mn8@2896_g N_VSS_Mn8@2896_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2897 N_OUT8_Mp8@2897_d N_OUT7_Mp8@2897_g N_VDD_Mp8@2897_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2896 N_OUT8_Mp8@2896_d N_OUT7_Mp8@2896_g N_VDD_Mp8@2896_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2895 N_OUT8_Mn8@2895_d N_OUT7_Mn8@2895_g N_VSS_Mn8@2895_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2894 N_OUT8_Mn8@2894_d N_OUT7_Mn8@2894_g N_VSS_Mn8@2894_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2895 N_OUT8_Mp8@2895_d N_OUT7_Mp8@2895_g N_VDD_Mp8@2895_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2894 N_OUT8_Mp8@2894_d N_OUT7_Mp8@2894_g N_VDD_Mp8@2894_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2893 N_OUT8_Mn8@2893_d N_OUT7_Mn8@2893_g N_VSS_Mn8@2893_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2892 N_OUT8_Mn8@2892_d N_OUT7_Mn8@2892_g N_VSS_Mn8@2892_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2893 N_OUT8_Mp8@2893_d N_OUT7_Mp8@2893_g N_VDD_Mp8@2893_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2892 N_OUT8_Mp8@2892_d N_OUT7_Mp8@2892_g N_VDD_Mp8@2892_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2891 N_OUT8_Mn8@2891_d N_OUT7_Mn8@2891_g N_VSS_Mn8@2891_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2890 N_OUT8_Mn8@2890_d N_OUT7_Mn8@2890_g N_VSS_Mn8@2890_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2891 N_OUT8_Mp8@2891_d N_OUT7_Mp8@2891_g N_VDD_Mp8@2891_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2890 N_OUT8_Mp8@2890_d N_OUT7_Mp8@2890_g N_VDD_Mp8@2890_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2889 N_OUT8_Mn8@2889_d N_OUT7_Mn8@2889_g N_VSS_Mn8@2889_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2888 N_OUT8_Mn8@2888_d N_OUT7_Mn8@2888_g N_VSS_Mn8@2888_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2889 N_OUT8_Mp8@2889_d N_OUT7_Mp8@2889_g N_VDD_Mp8@2889_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2888 N_OUT8_Mp8@2888_d N_OUT7_Mp8@2888_g N_VDD_Mp8@2888_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2887 N_OUT8_Mn8@2887_d N_OUT7_Mn8@2887_g N_VSS_Mn8@2887_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2886 N_OUT8_Mn8@2886_d N_OUT7_Mn8@2886_g N_VSS_Mn8@2886_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2887 N_OUT8_Mp8@2887_d N_OUT7_Mp8@2887_g N_VDD_Mp8@2887_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2886 N_OUT8_Mp8@2886_d N_OUT7_Mp8@2886_g N_VDD_Mp8@2886_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2885 N_OUT8_Mn8@2885_d N_OUT7_Mn8@2885_g N_VSS_Mn8@2885_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2884 N_OUT8_Mn8@2884_d N_OUT7_Mn8@2884_g N_VSS_Mn8@2884_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2885 N_OUT8_Mp8@2885_d N_OUT7_Mp8@2885_g N_VDD_Mp8@2885_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2884 N_OUT8_Mp8@2884_d N_OUT7_Mp8@2884_g N_VDD_Mp8@2884_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2883 N_OUT8_Mn8@2883_d N_OUT7_Mn8@2883_g N_VSS_Mn8@2883_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2882 N_OUT8_Mn8@2882_d N_OUT7_Mn8@2882_g N_VSS_Mn8@2882_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2883 N_OUT8_Mp8@2883_d N_OUT7_Mp8@2883_g N_VDD_Mp8@2883_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2882 N_OUT8_Mp8@2882_d N_OUT7_Mp8@2882_g N_VDD_Mp8@2882_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2881 N_OUT8_Mn8@2881_d N_OUT7_Mn8@2881_g N_VSS_Mn8@2881_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2880 N_OUT8_Mn8@2880_d N_OUT7_Mn8@2880_g N_VSS_Mn8@2880_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2881 N_OUT8_Mp8@2881_d N_OUT7_Mp8@2881_g N_VDD_Mp8@2881_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2880 N_OUT8_Mp8@2880_d N_OUT7_Mp8@2880_g N_VDD_Mp8@2880_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2879 N_OUT8_Mn8@2879_d N_OUT7_Mn8@2879_g N_VSS_Mn8@2879_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2878 N_OUT8_Mn8@2878_d N_OUT7_Mn8@2878_g N_VSS_Mn8@2878_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2879 N_OUT8_Mp8@2879_d N_OUT7_Mp8@2879_g N_VDD_Mp8@2879_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2878 N_OUT8_Mp8@2878_d N_OUT7_Mp8@2878_g N_VDD_Mp8@2878_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2877 N_OUT8_Mn8@2877_d N_OUT7_Mn8@2877_g N_VSS_Mn8@2877_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2876 N_OUT8_Mn8@2876_d N_OUT7_Mn8@2876_g N_VSS_Mn8@2876_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2877 N_OUT8_Mp8@2877_d N_OUT7_Mp8@2877_g N_VDD_Mp8@2877_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2876 N_OUT8_Mp8@2876_d N_OUT7_Mp8@2876_g N_VDD_Mp8@2876_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2875 N_OUT8_Mn8@2875_d N_OUT7_Mn8@2875_g N_VSS_Mn8@2875_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2874 N_OUT8_Mn8@2874_d N_OUT7_Mn8@2874_g N_VSS_Mn8@2874_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2875 N_OUT8_Mp8@2875_d N_OUT7_Mp8@2875_g N_VDD_Mp8@2875_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2874 N_OUT8_Mp8@2874_d N_OUT7_Mp8@2874_g N_VDD_Mp8@2874_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2873 N_OUT8_Mn8@2873_d N_OUT7_Mn8@2873_g N_VSS_Mn8@2873_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2872 N_OUT8_Mn8@2872_d N_OUT7_Mn8@2872_g N_VSS_Mn8@2872_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2873 N_OUT8_Mp8@2873_d N_OUT7_Mp8@2873_g N_VDD_Mp8@2873_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2872 N_OUT8_Mp8@2872_d N_OUT7_Mp8@2872_g N_VDD_Mp8@2872_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2871 N_OUT8_Mn8@2871_d N_OUT7_Mn8@2871_g N_VSS_Mn8@2871_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2870 N_OUT8_Mn8@2870_d N_OUT7_Mn8@2870_g N_VSS_Mn8@2870_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2871 N_OUT8_Mp8@2871_d N_OUT7_Mp8@2871_g N_VDD_Mp8@2871_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2870 N_OUT8_Mp8@2870_d N_OUT7_Mp8@2870_g N_VDD_Mp8@2870_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2869 N_OUT8_Mn8@2869_d N_OUT7_Mn8@2869_g N_VSS_Mn8@2869_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2868 N_OUT8_Mn8@2868_d N_OUT7_Mn8@2868_g N_VSS_Mn8@2868_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2869 N_OUT8_Mp8@2869_d N_OUT7_Mp8@2869_g N_VDD_Mp8@2869_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2868 N_OUT8_Mp8@2868_d N_OUT7_Mp8@2868_g N_VDD_Mp8@2868_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2867 N_OUT8_Mn8@2867_d N_OUT7_Mn8@2867_g N_VSS_Mn8@2867_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2866 N_OUT8_Mn8@2866_d N_OUT7_Mn8@2866_g N_VSS_Mn8@2866_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2867 N_OUT8_Mp8@2867_d N_OUT7_Mp8@2867_g N_VDD_Mp8@2867_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2866 N_OUT8_Mp8@2866_d N_OUT7_Mp8@2866_g N_VDD_Mp8@2866_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2865 N_OUT8_Mn8@2865_d N_OUT7_Mn8@2865_g N_VSS_Mn8@2865_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2864 N_OUT8_Mn8@2864_d N_OUT7_Mn8@2864_g N_VSS_Mn8@2864_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2865 N_OUT8_Mp8@2865_d N_OUT7_Mp8@2865_g N_VDD_Mp8@2865_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2864 N_OUT8_Mp8@2864_d N_OUT7_Mp8@2864_g N_VDD_Mp8@2864_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2863 N_OUT8_Mn8@2863_d N_OUT7_Mn8@2863_g N_VSS_Mn8@2863_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2862 N_OUT8_Mn8@2862_d N_OUT7_Mn8@2862_g N_VSS_Mn8@2862_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2863 N_OUT8_Mp8@2863_d N_OUT7_Mp8@2863_g N_VDD_Mp8@2863_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2862 N_OUT8_Mp8@2862_d N_OUT7_Mp8@2862_g N_VDD_Mp8@2862_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2861 N_OUT8_Mn8@2861_d N_OUT7_Mn8@2861_g N_VSS_Mn8@2861_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2860 N_OUT8_Mn8@2860_d N_OUT7_Mn8@2860_g N_VSS_Mn8@2860_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2861 N_OUT8_Mp8@2861_d N_OUT7_Mp8@2861_g N_VDD_Mp8@2861_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2860 N_OUT8_Mp8@2860_d N_OUT7_Mp8@2860_g N_VDD_Mp8@2860_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2859 N_OUT8_Mn8@2859_d N_OUT7_Mn8@2859_g N_VSS_Mn8@2859_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2858 N_OUT8_Mn8@2858_d N_OUT7_Mn8@2858_g N_VSS_Mn8@2858_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2859 N_OUT8_Mp8@2859_d N_OUT7_Mp8@2859_g N_VDD_Mp8@2859_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2858 N_OUT8_Mp8@2858_d N_OUT7_Mp8@2858_g N_VDD_Mp8@2858_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2857 N_OUT8_Mn8@2857_d N_OUT7_Mn8@2857_g N_VSS_Mn8@2857_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2856 N_OUT8_Mn8@2856_d N_OUT7_Mn8@2856_g N_VSS_Mn8@2856_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2857 N_OUT8_Mp8@2857_d N_OUT7_Mp8@2857_g N_VDD_Mp8@2857_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2856 N_OUT8_Mp8@2856_d N_OUT7_Mp8@2856_g N_VDD_Mp8@2856_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2855 N_OUT8_Mn8@2855_d N_OUT7_Mn8@2855_g N_VSS_Mn8@2855_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2854 N_OUT8_Mn8@2854_d N_OUT7_Mn8@2854_g N_VSS_Mn8@2854_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2855 N_OUT8_Mp8@2855_d N_OUT7_Mp8@2855_g N_VDD_Mp8@2855_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2854 N_OUT8_Mp8@2854_d N_OUT7_Mp8@2854_g N_VDD_Mp8@2854_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2853 N_OUT8_Mn8@2853_d N_OUT7_Mn8@2853_g N_VSS_Mn8@2853_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2852 N_OUT8_Mn8@2852_d N_OUT7_Mn8@2852_g N_VSS_Mn8@2852_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2853 N_OUT8_Mp8@2853_d N_OUT7_Mp8@2853_g N_VDD_Mp8@2853_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2852 N_OUT8_Mp8@2852_d N_OUT7_Mp8@2852_g N_VDD_Mp8@2852_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2851 N_OUT8_Mn8@2851_d N_OUT7_Mn8@2851_g N_VSS_Mn8@2851_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2850 N_OUT8_Mn8@2850_d N_OUT7_Mn8@2850_g N_VSS_Mn8@2850_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2851 N_OUT8_Mp8@2851_d N_OUT7_Mp8@2851_g N_VDD_Mp8@2851_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2850 N_OUT8_Mp8@2850_d N_OUT7_Mp8@2850_g N_VDD_Mp8@2850_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2849 N_OUT8_Mn8@2849_d N_OUT7_Mn8@2849_g N_VSS_Mn8@2849_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2848 N_OUT8_Mn8@2848_d N_OUT7_Mn8@2848_g N_VSS_Mn8@2848_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2849 N_OUT8_Mp8@2849_d N_OUT7_Mp8@2849_g N_VDD_Mp8@2849_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2848 N_OUT8_Mp8@2848_d N_OUT7_Mp8@2848_g N_VDD_Mp8@2848_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2847 N_OUT8_Mn8@2847_d N_OUT7_Mn8@2847_g N_VSS_Mn8@2847_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2846 N_OUT8_Mn8@2846_d N_OUT7_Mn8@2846_g N_VSS_Mn8@2846_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2847 N_OUT8_Mp8@2847_d N_OUT7_Mp8@2847_g N_VDD_Mp8@2847_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2846 N_OUT8_Mp8@2846_d N_OUT7_Mp8@2846_g N_VDD_Mp8@2846_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2845 N_OUT8_Mn8@2845_d N_OUT7_Mn8@2845_g N_VSS_Mn8@2845_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2844 N_OUT8_Mn8@2844_d N_OUT7_Mn8@2844_g N_VSS_Mn8@2844_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2845 N_OUT8_Mp8@2845_d N_OUT7_Mp8@2845_g N_VDD_Mp8@2845_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2844 N_OUT8_Mp8@2844_d N_OUT7_Mp8@2844_g N_VDD_Mp8@2844_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2843 N_OUT8_Mn8@2843_d N_OUT7_Mn8@2843_g N_VSS_Mn8@2843_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2842 N_OUT8_Mn8@2842_d N_OUT7_Mn8@2842_g N_VSS_Mn8@2842_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2843 N_OUT8_Mp8@2843_d N_OUT7_Mp8@2843_g N_VDD_Mp8@2843_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2842 N_OUT8_Mp8@2842_d N_OUT7_Mp8@2842_g N_VDD_Mp8@2842_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2841 N_OUT8_Mn8@2841_d N_OUT7_Mn8@2841_g N_VSS_Mn8@2841_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2840 N_OUT8_Mn8@2840_d N_OUT7_Mn8@2840_g N_VSS_Mn8@2840_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2841 N_OUT8_Mp8@2841_d N_OUT7_Mp8@2841_g N_VDD_Mp8@2841_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2840 N_OUT8_Mp8@2840_d N_OUT7_Mp8@2840_g N_VDD_Mp8@2840_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2839 N_OUT8_Mn8@2839_d N_OUT7_Mn8@2839_g N_VSS_Mn8@2839_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2838 N_OUT8_Mn8@2838_d N_OUT7_Mn8@2838_g N_VSS_Mn8@2838_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2839 N_OUT8_Mp8@2839_d N_OUT7_Mp8@2839_g N_VDD_Mp8@2839_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2838 N_OUT8_Mp8@2838_d N_OUT7_Mp8@2838_g N_VDD_Mp8@2838_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2837 N_OUT8_Mn8@2837_d N_OUT7_Mn8@2837_g N_VSS_Mn8@2837_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2836 N_OUT8_Mn8@2836_d N_OUT7_Mn8@2836_g N_VSS_Mn8@2836_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2837 N_OUT8_Mp8@2837_d N_OUT7_Mp8@2837_g N_VDD_Mp8@2837_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2836 N_OUT8_Mp8@2836_d N_OUT7_Mp8@2836_g N_VDD_Mp8@2836_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2835 N_OUT8_Mn8@2835_d N_OUT7_Mn8@2835_g N_VSS_Mn8@2835_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2834 N_OUT8_Mn8@2834_d N_OUT7_Mn8@2834_g N_VSS_Mn8@2834_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2835 N_OUT8_Mp8@2835_d N_OUT7_Mp8@2835_g N_VDD_Mp8@2835_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2834 N_OUT8_Mp8@2834_d N_OUT7_Mp8@2834_g N_VDD_Mp8@2834_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2833 N_OUT8_Mn8@2833_d N_OUT7_Mn8@2833_g N_VSS_Mn8@2833_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2832 N_OUT8_Mn8@2832_d N_OUT7_Mn8@2832_g N_VSS_Mn8@2832_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2833 N_OUT8_Mp8@2833_d N_OUT7_Mp8@2833_g N_VDD_Mp8@2833_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2832 N_OUT8_Mp8@2832_d N_OUT7_Mp8@2832_g N_VDD_Mp8@2832_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2831 N_OUT8_Mn8@2831_d N_OUT7_Mn8@2831_g N_VSS_Mn8@2831_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2830 N_OUT8_Mn8@2830_d N_OUT7_Mn8@2830_g N_VSS_Mn8@2830_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2831 N_OUT8_Mp8@2831_d N_OUT7_Mp8@2831_g N_VDD_Mp8@2831_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2830 N_OUT8_Mp8@2830_d N_OUT7_Mp8@2830_g N_VDD_Mp8@2830_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2829 N_OUT8_Mn8@2829_d N_OUT7_Mn8@2829_g N_VSS_Mn8@2829_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2828 N_OUT8_Mn8@2828_d N_OUT7_Mn8@2828_g N_VSS_Mn8@2828_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2829 N_OUT8_Mp8@2829_d N_OUT7_Mp8@2829_g N_VDD_Mp8@2829_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2828 N_OUT8_Mp8@2828_d N_OUT7_Mp8@2828_g N_VDD_Mp8@2828_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2827 N_OUT8_Mn8@2827_d N_OUT7_Mn8@2827_g N_VSS_Mn8@2827_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2826 N_OUT8_Mn8@2826_d N_OUT7_Mn8@2826_g N_VSS_Mn8@2826_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2827 N_OUT8_Mp8@2827_d N_OUT7_Mp8@2827_g N_VDD_Mp8@2827_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2826 N_OUT8_Mp8@2826_d N_OUT7_Mp8@2826_g N_VDD_Mp8@2826_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2825 N_OUT8_Mn8@2825_d N_OUT7_Mn8@2825_g N_VSS_Mn8@2825_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2824 N_OUT8_Mn8@2824_d N_OUT7_Mn8@2824_g N_VSS_Mn8@2824_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2825 N_OUT8_Mp8@2825_d N_OUT7_Mp8@2825_g N_VDD_Mp8@2825_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2824 N_OUT8_Mp8@2824_d N_OUT7_Mp8@2824_g N_VDD_Mp8@2824_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2823 N_OUT8_Mn8@2823_d N_OUT7_Mn8@2823_g N_VSS_Mn8@2823_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2822 N_OUT8_Mn8@2822_d N_OUT7_Mn8@2822_g N_VSS_Mn8@2822_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2823 N_OUT8_Mp8@2823_d N_OUT7_Mp8@2823_g N_VDD_Mp8@2823_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2822 N_OUT8_Mp8@2822_d N_OUT7_Mp8@2822_g N_VDD_Mp8@2822_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2821 N_OUT8_Mn8@2821_d N_OUT7_Mn8@2821_g N_VSS_Mn8@2821_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2820 N_OUT8_Mn8@2820_d N_OUT7_Mn8@2820_g N_VSS_Mn8@2820_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2821 N_OUT8_Mp8@2821_d N_OUT7_Mp8@2821_g N_VDD_Mp8@2821_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2820 N_OUT8_Mp8@2820_d N_OUT7_Mp8@2820_g N_VDD_Mp8@2820_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2819 N_OUT8_Mn8@2819_d N_OUT7_Mn8@2819_g N_VSS_Mn8@2819_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2818 N_OUT8_Mn8@2818_d N_OUT7_Mn8@2818_g N_VSS_Mn8@2818_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2819 N_OUT8_Mp8@2819_d N_OUT7_Mp8@2819_g N_VDD_Mp8@2819_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2818 N_OUT8_Mp8@2818_d N_OUT7_Mp8@2818_g N_VDD_Mp8@2818_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2817 N_OUT8_Mn8@2817_d N_OUT7_Mn8@2817_g N_VSS_Mn8@2817_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2816 N_OUT8_Mn8@2816_d N_OUT7_Mn8@2816_g N_VSS_Mn8@2816_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2817 N_OUT8_Mp8@2817_d N_OUT7_Mp8@2817_g N_VDD_Mp8@2817_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2816 N_OUT8_Mp8@2816_d N_OUT7_Mp8@2816_g N_VDD_Mp8@2816_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2815 N_OUT8_Mn8@2815_d N_OUT7_Mn8@2815_g N_VSS_Mn8@2815_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2814 N_OUT8_Mn8@2814_d N_OUT7_Mn8@2814_g N_VSS_Mn8@2814_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2815 N_OUT8_Mp8@2815_d N_OUT7_Mp8@2815_g N_VDD_Mp8@2815_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2814 N_OUT8_Mp8@2814_d N_OUT7_Mp8@2814_g N_VDD_Mp8@2814_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2813 N_OUT8_Mn8@2813_d N_OUT7_Mn8@2813_g N_VSS_Mn8@2813_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2812 N_OUT8_Mn8@2812_d N_OUT7_Mn8@2812_g N_VSS_Mn8@2812_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2813 N_OUT8_Mp8@2813_d N_OUT7_Mp8@2813_g N_VDD_Mp8@2813_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2812 N_OUT8_Mp8@2812_d N_OUT7_Mp8@2812_g N_VDD_Mp8@2812_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2811 N_OUT8_Mn8@2811_d N_OUT7_Mn8@2811_g N_VSS_Mn8@2811_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2810 N_OUT8_Mn8@2810_d N_OUT7_Mn8@2810_g N_VSS_Mn8@2810_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2811 N_OUT8_Mp8@2811_d N_OUT7_Mp8@2811_g N_VDD_Mp8@2811_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2810 N_OUT8_Mp8@2810_d N_OUT7_Mp8@2810_g N_VDD_Mp8@2810_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2809 N_OUT8_Mn8@2809_d N_OUT7_Mn8@2809_g N_VSS_Mn8@2809_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2808 N_OUT8_Mn8@2808_d N_OUT7_Mn8@2808_g N_VSS_Mn8@2808_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2809 N_OUT8_Mp8@2809_d N_OUT7_Mp8@2809_g N_VDD_Mp8@2809_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2808 N_OUT8_Mp8@2808_d N_OUT7_Mp8@2808_g N_VDD_Mp8@2808_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2807 N_OUT8_Mn8@2807_d N_OUT7_Mn8@2807_g N_VSS_Mn8@2807_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2806 N_OUT8_Mn8@2806_d N_OUT7_Mn8@2806_g N_VSS_Mn8@2806_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2807 N_OUT8_Mp8@2807_d N_OUT7_Mp8@2807_g N_VDD_Mp8@2807_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2806 N_OUT8_Mp8@2806_d N_OUT7_Mp8@2806_g N_VDD_Mp8@2806_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2805 N_OUT8_Mn8@2805_d N_OUT7_Mn8@2805_g N_VSS_Mn8@2805_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2804 N_OUT8_Mn8@2804_d N_OUT7_Mn8@2804_g N_VSS_Mn8@2804_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2805 N_OUT8_Mp8@2805_d N_OUT7_Mp8@2805_g N_VDD_Mp8@2805_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2804 N_OUT8_Mp8@2804_d N_OUT7_Mp8@2804_g N_VDD_Mp8@2804_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2803 N_OUT8_Mn8@2803_d N_OUT7_Mn8@2803_g N_VSS_Mn8@2803_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2802 N_OUT8_Mn8@2802_d N_OUT7_Mn8@2802_g N_VSS_Mn8@2802_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2803 N_OUT8_Mp8@2803_d N_OUT7_Mp8@2803_g N_VDD_Mp8@2803_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2802 N_OUT8_Mp8@2802_d N_OUT7_Mp8@2802_g N_VDD_Mp8@2802_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2801 N_OUT8_Mn8@2801_d N_OUT7_Mn8@2801_g N_VSS_Mn8@2801_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2800 N_OUT8_Mn8@2800_d N_OUT7_Mn8@2800_g N_VSS_Mn8@2800_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2801 N_OUT8_Mp8@2801_d N_OUT7_Mp8@2801_g N_VDD_Mp8@2801_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2800 N_OUT8_Mp8@2800_d N_OUT7_Mp8@2800_g N_VDD_Mp8@2800_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2799 N_OUT8_Mn8@2799_d N_OUT7_Mn8@2799_g N_VSS_Mn8@2799_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2798 N_OUT8_Mn8@2798_d N_OUT7_Mn8@2798_g N_VSS_Mn8@2798_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2799 N_OUT8_Mp8@2799_d N_OUT7_Mp8@2799_g N_VDD_Mp8@2799_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2798 N_OUT8_Mp8@2798_d N_OUT7_Mp8@2798_g N_VDD_Mp8@2798_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2797 N_OUT8_Mn8@2797_d N_OUT7_Mn8@2797_g N_VSS_Mn8@2797_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2796 N_OUT8_Mn8@2796_d N_OUT7_Mn8@2796_g N_VSS_Mn8@2796_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2797 N_OUT8_Mp8@2797_d N_OUT7_Mp8@2797_g N_VDD_Mp8@2797_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2796 N_OUT8_Mp8@2796_d N_OUT7_Mp8@2796_g N_VDD_Mp8@2796_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2795 N_OUT8_Mn8@2795_d N_OUT7_Mn8@2795_g N_VSS_Mn8@2795_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2794 N_OUT8_Mn8@2794_d N_OUT7_Mn8@2794_g N_VSS_Mn8@2794_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2795 N_OUT8_Mp8@2795_d N_OUT7_Mp8@2795_g N_VDD_Mp8@2795_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2794 N_OUT8_Mp8@2794_d N_OUT7_Mp8@2794_g N_VDD_Mp8@2794_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2793 N_OUT8_Mn8@2793_d N_OUT7_Mn8@2793_g N_VSS_Mn8@2793_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2792 N_OUT8_Mn8@2792_d N_OUT7_Mn8@2792_g N_VSS_Mn8@2792_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2793 N_OUT8_Mp8@2793_d N_OUT7_Mp8@2793_g N_VDD_Mp8@2793_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2792 N_OUT8_Mp8@2792_d N_OUT7_Mp8@2792_g N_VDD_Mp8@2792_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2791 N_OUT8_Mn8@2791_d N_OUT7_Mn8@2791_g N_VSS_Mn8@2791_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2790 N_OUT8_Mn8@2790_d N_OUT7_Mn8@2790_g N_VSS_Mn8@2790_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2791 N_OUT8_Mp8@2791_d N_OUT7_Mp8@2791_g N_VDD_Mp8@2791_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2790 N_OUT8_Mp8@2790_d N_OUT7_Mp8@2790_g N_VDD_Mp8@2790_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2789 N_OUT8_Mn8@2789_d N_OUT7_Mn8@2789_g N_VSS_Mn8@2789_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2788 N_OUT8_Mn8@2788_d N_OUT7_Mn8@2788_g N_VSS_Mn8@2788_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2789 N_OUT8_Mp8@2789_d N_OUT7_Mp8@2789_g N_VDD_Mp8@2789_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2788 N_OUT8_Mp8@2788_d N_OUT7_Mp8@2788_g N_VDD_Mp8@2788_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2787 N_OUT8_Mn8@2787_d N_OUT7_Mn8@2787_g N_VSS_Mn8@2787_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2786 N_OUT8_Mn8@2786_d N_OUT7_Mn8@2786_g N_VSS_Mn8@2786_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2787 N_OUT8_Mp8@2787_d N_OUT7_Mp8@2787_g N_VDD_Mp8@2787_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2786 N_OUT8_Mp8@2786_d N_OUT7_Mp8@2786_g N_VDD_Mp8@2786_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2785 N_OUT8_Mn8@2785_d N_OUT7_Mn8@2785_g N_VSS_Mn8@2785_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2784 N_OUT8_Mn8@2784_d N_OUT7_Mn8@2784_g N_VSS_Mn8@2784_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2785 N_OUT8_Mp8@2785_d N_OUT7_Mp8@2785_g N_VDD_Mp8@2785_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2784 N_OUT8_Mp8@2784_d N_OUT7_Mp8@2784_g N_VDD_Mp8@2784_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2783 N_OUT8_Mn8@2783_d N_OUT7_Mn8@2783_g N_VSS_Mn8@2783_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2782 N_OUT8_Mn8@2782_d N_OUT7_Mn8@2782_g N_VSS_Mn8@2782_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2783 N_OUT8_Mp8@2783_d N_OUT7_Mp8@2783_g N_VDD_Mp8@2783_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2782 N_OUT8_Mp8@2782_d N_OUT7_Mp8@2782_g N_VDD_Mp8@2782_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2781 N_OUT8_Mn8@2781_d N_OUT7_Mn8@2781_g N_VSS_Mn8@2781_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2780 N_OUT8_Mn8@2780_d N_OUT7_Mn8@2780_g N_VSS_Mn8@2780_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2781 N_OUT8_Mp8@2781_d N_OUT7_Mp8@2781_g N_VDD_Mp8@2781_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2780 N_OUT8_Mp8@2780_d N_OUT7_Mp8@2780_g N_VDD_Mp8@2780_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2779 N_OUT8_Mn8@2779_d N_OUT7_Mn8@2779_g N_VSS_Mn8@2779_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2778 N_OUT8_Mn8@2778_d N_OUT7_Mn8@2778_g N_VSS_Mn8@2778_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2779 N_OUT8_Mp8@2779_d N_OUT7_Mp8@2779_g N_VDD_Mp8@2779_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2778 N_OUT8_Mp8@2778_d N_OUT7_Mp8@2778_g N_VDD_Mp8@2778_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2777 N_OUT8_Mn8@2777_d N_OUT7_Mn8@2777_g N_VSS_Mn8@2777_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2776 N_OUT8_Mn8@2776_d N_OUT7_Mn8@2776_g N_VSS_Mn8@2776_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2777 N_OUT8_Mp8@2777_d N_OUT7_Mp8@2777_g N_VDD_Mp8@2777_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2776 N_OUT8_Mp8@2776_d N_OUT7_Mp8@2776_g N_VDD_Mp8@2776_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2775 N_OUT8_Mn8@2775_d N_OUT7_Mn8@2775_g N_VSS_Mn8@2775_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2774 N_OUT8_Mn8@2774_d N_OUT7_Mn8@2774_g N_VSS_Mn8@2774_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2775 N_OUT8_Mp8@2775_d N_OUT7_Mp8@2775_g N_VDD_Mp8@2775_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2774 N_OUT8_Mp8@2774_d N_OUT7_Mp8@2774_g N_VDD_Mp8@2774_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2773 N_OUT8_Mn8@2773_d N_OUT7_Mn8@2773_g N_VSS_Mn8@2773_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2772 N_OUT8_Mn8@2772_d N_OUT7_Mn8@2772_g N_VSS_Mn8@2772_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2773 N_OUT8_Mp8@2773_d N_OUT7_Mp8@2773_g N_VDD_Mp8@2773_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2772 N_OUT8_Mp8@2772_d N_OUT7_Mp8@2772_g N_VDD_Mp8@2772_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2771 N_OUT8_Mn8@2771_d N_OUT7_Mn8@2771_g N_VSS_Mn8@2771_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2770 N_OUT8_Mn8@2770_d N_OUT7_Mn8@2770_g N_VSS_Mn8@2770_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2771 N_OUT8_Mp8@2771_d N_OUT7_Mp8@2771_g N_VDD_Mp8@2771_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2770 N_OUT8_Mp8@2770_d N_OUT7_Mp8@2770_g N_VDD_Mp8@2770_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2769 N_OUT8_Mn8@2769_d N_OUT7_Mn8@2769_g N_VSS_Mn8@2769_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2768 N_OUT8_Mn8@2768_d N_OUT7_Mn8@2768_g N_VSS_Mn8@2768_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2769 N_OUT8_Mp8@2769_d N_OUT7_Mp8@2769_g N_VDD_Mp8@2769_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2768 N_OUT8_Mp8@2768_d N_OUT7_Mp8@2768_g N_VDD_Mp8@2768_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2767 N_OUT8_Mn8@2767_d N_OUT7_Mn8@2767_g N_VSS_Mn8@2767_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2766 N_OUT8_Mn8@2766_d N_OUT7_Mn8@2766_g N_VSS_Mn8@2766_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2767 N_OUT8_Mp8@2767_d N_OUT7_Mp8@2767_g N_VDD_Mp8@2767_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2766 N_OUT8_Mp8@2766_d N_OUT7_Mp8@2766_g N_VDD_Mp8@2766_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2765 N_OUT8_Mn8@2765_d N_OUT7_Mn8@2765_g N_VSS_Mn8@2765_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2764 N_OUT8_Mn8@2764_d N_OUT7_Mn8@2764_g N_VSS_Mn8@2764_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2765 N_OUT8_Mp8@2765_d N_OUT7_Mp8@2765_g N_VDD_Mp8@2765_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2764 N_OUT8_Mp8@2764_d N_OUT7_Mp8@2764_g N_VDD_Mp8@2764_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2763 N_OUT8_Mn8@2763_d N_OUT7_Mn8@2763_g N_VSS_Mn8@2763_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2762 N_OUT8_Mn8@2762_d N_OUT7_Mn8@2762_g N_VSS_Mn8@2762_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2763 N_OUT8_Mp8@2763_d N_OUT7_Mp8@2763_g N_VDD_Mp8@2763_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2762 N_OUT8_Mp8@2762_d N_OUT7_Mp8@2762_g N_VDD_Mp8@2762_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2761 N_OUT8_Mn8@2761_d N_OUT7_Mn8@2761_g N_VSS_Mn8@2761_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2760 N_OUT8_Mn8@2760_d N_OUT7_Mn8@2760_g N_VSS_Mn8@2760_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2761 N_OUT8_Mp8@2761_d N_OUT7_Mp8@2761_g N_VDD_Mp8@2761_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2760 N_OUT8_Mp8@2760_d N_OUT7_Mp8@2760_g N_VDD_Mp8@2760_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2759 N_OUT8_Mn8@2759_d N_OUT7_Mn8@2759_g N_VSS_Mn8@2759_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2758 N_OUT8_Mn8@2758_d N_OUT7_Mn8@2758_g N_VSS_Mn8@2758_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2759 N_OUT8_Mp8@2759_d N_OUT7_Mp8@2759_g N_VDD_Mp8@2759_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2758 N_OUT8_Mp8@2758_d N_OUT7_Mp8@2758_g N_VDD_Mp8@2758_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2757 N_OUT8_Mn8@2757_d N_OUT7_Mn8@2757_g N_VSS_Mn8@2757_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2756 N_OUT8_Mn8@2756_d N_OUT7_Mn8@2756_g N_VSS_Mn8@2756_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2757 N_OUT8_Mp8@2757_d N_OUT7_Mp8@2757_g N_VDD_Mp8@2757_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2756 N_OUT8_Mp8@2756_d N_OUT7_Mp8@2756_g N_VDD_Mp8@2756_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2755 N_OUT8_Mn8@2755_d N_OUT7_Mn8@2755_g N_VSS_Mn8@2755_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2754 N_OUT8_Mn8@2754_d N_OUT7_Mn8@2754_g N_VSS_Mn8@2754_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2755 N_OUT8_Mp8@2755_d N_OUT7_Mp8@2755_g N_VDD_Mp8@2755_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2754 N_OUT8_Mp8@2754_d N_OUT7_Mp8@2754_g N_VDD_Mp8@2754_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2753 N_OUT8_Mn8@2753_d N_OUT7_Mn8@2753_g N_VSS_Mn8@2753_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2752 N_OUT8_Mn8@2752_d N_OUT7_Mn8@2752_g N_VSS_Mn8@2752_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2753 N_OUT8_Mp8@2753_d N_OUT7_Mp8@2753_g N_VDD_Mp8@2753_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2752 N_OUT8_Mp8@2752_d N_OUT7_Mp8@2752_g N_VDD_Mp8@2752_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2751 N_OUT8_Mn8@2751_d N_OUT7_Mn8@2751_g N_VSS_Mn8@2751_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2750 N_OUT8_Mn8@2750_d N_OUT7_Mn8@2750_g N_VSS_Mn8@2750_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2751 N_OUT8_Mp8@2751_d N_OUT7_Mp8@2751_g N_VDD_Mp8@2751_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2750 N_OUT8_Mp8@2750_d N_OUT7_Mp8@2750_g N_VDD_Mp8@2750_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2749 N_OUT8_Mn8@2749_d N_OUT7_Mn8@2749_g N_VSS_Mn8@2749_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2748 N_OUT8_Mn8@2748_d N_OUT7_Mn8@2748_g N_VSS_Mn8@2748_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2749 N_OUT8_Mp8@2749_d N_OUT7_Mp8@2749_g N_VDD_Mp8@2749_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2748 N_OUT8_Mp8@2748_d N_OUT7_Mp8@2748_g N_VDD_Mp8@2748_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2747 N_OUT8_Mn8@2747_d N_OUT7_Mn8@2747_g N_VSS_Mn8@2747_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2746 N_OUT8_Mn8@2746_d N_OUT7_Mn8@2746_g N_VSS_Mn8@2746_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2747 N_OUT8_Mp8@2747_d N_OUT7_Mp8@2747_g N_VDD_Mp8@2747_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2746 N_OUT8_Mp8@2746_d N_OUT7_Mp8@2746_g N_VDD_Mp8@2746_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2745 N_OUT8_Mn8@2745_d N_OUT7_Mn8@2745_g N_VSS_Mn8@2745_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2744 N_OUT8_Mn8@2744_d N_OUT7_Mn8@2744_g N_VSS_Mn8@2744_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2745 N_OUT8_Mp8@2745_d N_OUT7_Mp8@2745_g N_VDD_Mp8@2745_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2744 N_OUT8_Mp8@2744_d N_OUT7_Mp8@2744_g N_VDD_Mp8@2744_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2743 N_OUT8_Mn8@2743_d N_OUT7_Mn8@2743_g N_VSS_Mn8@2743_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2742 N_OUT8_Mn8@2742_d N_OUT7_Mn8@2742_g N_VSS_Mn8@2742_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2743 N_OUT8_Mp8@2743_d N_OUT7_Mp8@2743_g N_VDD_Mp8@2743_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2742 N_OUT8_Mp8@2742_d N_OUT7_Mp8@2742_g N_VDD_Mp8@2742_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2741 N_OUT8_Mn8@2741_d N_OUT7_Mn8@2741_g N_VSS_Mn8@2741_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2740 N_OUT8_Mn8@2740_d N_OUT7_Mn8@2740_g N_VSS_Mn8@2740_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2741 N_OUT8_Mp8@2741_d N_OUT7_Mp8@2741_g N_VDD_Mp8@2741_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2740 N_OUT8_Mp8@2740_d N_OUT7_Mp8@2740_g N_VDD_Mp8@2740_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2739 N_OUT8_Mn8@2739_d N_OUT7_Mn8@2739_g N_VSS_Mn8@2739_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2738 N_OUT8_Mn8@2738_d N_OUT7_Mn8@2738_g N_VSS_Mn8@2738_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2739 N_OUT8_Mp8@2739_d N_OUT7_Mp8@2739_g N_VDD_Mp8@2739_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2738 N_OUT8_Mp8@2738_d N_OUT7_Mp8@2738_g N_VDD_Mp8@2738_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2737 N_OUT8_Mn8@2737_d N_OUT7_Mn8@2737_g N_VSS_Mn8@2737_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2736 N_OUT8_Mn8@2736_d N_OUT7_Mn8@2736_g N_VSS_Mn8@2736_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2737 N_OUT8_Mp8@2737_d N_OUT7_Mp8@2737_g N_VDD_Mp8@2737_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2736 N_OUT8_Mp8@2736_d N_OUT7_Mp8@2736_g N_VDD_Mp8@2736_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2735 N_OUT8_Mn8@2735_d N_OUT7_Mn8@2735_g N_VSS_Mn8@2735_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2734 N_OUT8_Mn8@2734_d N_OUT7_Mn8@2734_g N_VSS_Mn8@2734_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2735 N_OUT8_Mp8@2735_d N_OUT7_Mp8@2735_g N_VDD_Mp8@2735_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2734 N_OUT8_Mp8@2734_d N_OUT7_Mp8@2734_g N_VDD_Mp8@2734_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2733 N_OUT8_Mn8@2733_d N_OUT7_Mn8@2733_g N_VSS_Mn8@2733_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2732 N_OUT8_Mn8@2732_d N_OUT7_Mn8@2732_g N_VSS_Mn8@2732_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2733 N_OUT8_Mp8@2733_d N_OUT7_Mp8@2733_g N_VDD_Mp8@2733_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2732 N_OUT8_Mp8@2732_d N_OUT7_Mp8@2732_g N_VDD_Mp8@2732_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2731 N_OUT8_Mn8@2731_d N_OUT7_Mn8@2731_g N_VSS_Mn8@2731_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2730 N_OUT8_Mn8@2730_d N_OUT7_Mn8@2730_g N_VSS_Mn8@2730_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2731 N_OUT8_Mp8@2731_d N_OUT7_Mp8@2731_g N_VDD_Mp8@2731_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2730 N_OUT8_Mp8@2730_d N_OUT7_Mp8@2730_g N_VDD_Mp8@2730_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2729 N_OUT8_Mn8@2729_d N_OUT7_Mn8@2729_g N_VSS_Mn8@2729_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2728 N_OUT8_Mn8@2728_d N_OUT7_Mn8@2728_g N_VSS_Mn8@2728_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2729 N_OUT8_Mp8@2729_d N_OUT7_Mp8@2729_g N_VDD_Mp8@2729_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2728 N_OUT8_Mp8@2728_d N_OUT7_Mp8@2728_g N_VDD_Mp8@2728_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2727 N_OUT8_Mn8@2727_d N_OUT7_Mn8@2727_g N_VSS_Mn8@2727_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2726 N_OUT8_Mn8@2726_d N_OUT7_Mn8@2726_g N_VSS_Mn8@2726_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2727 N_OUT8_Mp8@2727_d N_OUT7_Mp8@2727_g N_VDD_Mp8@2727_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2726 N_OUT8_Mp8@2726_d N_OUT7_Mp8@2726_g N_VDD_Mp8@2726_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2725 N_OUT8_Mn8@2725_d N_OUT7_Mn8@2725_g N_VSS_Mn8@2725_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2724 N_OUT8_Mn8@2724_d N_OUT7_Mn8@2724_g N_VSS_Mn8@2724_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2725 N_OUT8_Mp8@2725_d N_OUT7_Mp8@2725_g N_VDD_Mp8@2725_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2724 N_OUT8_Mp8@2724_d N_OUT7_Mp8@2724_g N_VDD_Mp8@2724_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2723 N_OUT8_Mn8@2723_d N_OUT7_Mn8@2723_g N_VSS_Mn8@2723_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2722 N_OUT8_Mn8@2722_d N_OUT7_Mn8@2722_g N_VSS_Mn8@2722_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2723 N_OUT8_Mp8@2723_d N_OUT7_Mp8@2723_g N_VDD_Mp8@2723_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2722 N_OUT8_Mp8@2722_d N_OUT7_Mp8@2722_g N_VDD_Mp8@2722_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2721 N_OUT8_Mn8@2721_d N_OUT7_Mn8@2721_g N_VSS_Mn8@2721_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2720 N_OUT8_Mn8@2720_d N_OUT7_Mn8@2720_g N_VSS_Mn8@2720_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2721 N_OUT8_Mp8@2721_d N_OUT7_Mp8@2721_g N_VDD_Mp8@2721_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2720 N_OUT8_Mp8@2720_d N_OUT7_Mp8@2720_g N_VDD_Mp8@2720_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2719 N_OUT8_Mn8@2719_d N_OUT7_Mn8@2719_g N_VSS_Mn8@2719_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2718 N_OUT8_Mn8@2718_d N_OUT7_Mn8@2718_g N_VSS_Mn8@2718_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2719 N_OUT8_Mp8@2719_d N_OUT7_Mp8@2719_g N_VDD_Mp8@2719_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2718 N_OUT8_Mp8@2718_d N_OUT7_Mp8@2718_g N_VDD_Mp8@2718_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2717 N_OUT8_Mn8@2717_d N_OUT7_Mn8@2717_g N_VSS_Mn8@2717_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2716 N_OUT8_Mn8@2716_d N_OUT7_Mn8@2716_g N_VSS_Mn8@2716_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2717 N_OUT8_Mp8@2717_d N_OUT7_Mp8@2717_g N_VDD_Mp8@2717_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2716 N_OUT8_Mp8@2716_d N_OUT7_Mp8@2716_g N_VDD_Mp8@2716_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2715 N_OUT8_Mn8@2715_d N_OUT7_Mn8@2715_g N_VSS_Mn8@2715_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2714 N_OUT8_Mn8@2714_d N_OUT7_Mn8@2714_g N_VSS_Mn8@2714_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2715 N_OUT8_Mp8@2715_d N_OUT7_Mp8@2715_g N_VDD_Mp8@2715_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2714 N_OUT8_Mp8@2714_d N_OUT7_Mp8@2714_g N_VDD_Mp8@2714_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2713 N_OUT8_Mn8@2713_d N_OUT7_Mn8@2713_g N_VSS_Mn8@2713_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2712 N_OUT8_Mn8@2712_d N_OUT7_Mn8@2712_g N_VSS_Mn8@2712_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2713 N_OUT8_Mp8@2713_d N_OUT7_Mp8@2713_g N_VDD_Mp8@2713_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2712 N_OUT8_Mp8@2712_d N_OUT7_Mp8@2712_g N_VDD_Mp8@2712_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2711 N_OUT8_Mn8@2711_d N_OUT7_Mn8@2711_g N_VSS_Mn8@2711_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2710 N_OUT8_Mn8@2710_d N_OUT7_Mn8@2710_g N_VSS_Mn8@2710_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2711 N_OUT8_Mp8@2711_d N_OUT7_Mp8@2711_g N_VDD_Mp8@2711_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2710 N_OUT8_Mp8@2710_d N_OUT7_Mp8@2710_g N_VDD_Mp8@2710_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2709 N_OUT8_Mn8@2709_d N_OUT7_Mn8@2709_g N_VSS_Mn8@2709_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2708 N_OUT8_Mn8@2708_d N_OUT7_Mn8@2708_g N_VSS_Mn8@2708_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2709 N_OUT8_Mp8@2709_d N_OUT7_Mp8@2709_g N_VDD_Mp8@2709_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2708 N_OUT8_Mp8@2708_d N_OUT7_Mp8@2708_g N_VDD_Mp8@2708_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2707 N_OUT8_Mn8@2707_d N_OUT7_Mn8@2707_g N_VSS_Mn8@2707_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2706 N_OUT8_Mn8@2706_d N_OUT7_Mn8@2706_g N_VSS_Mn8@2706_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2707 N_OUT8_Mp8@2707_d N_OUT7_Mp8@2707_g N_VDD_Mp8@2707_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2706 N_OUT8_Mp8@2706_d N_OUT7_Mp8@2706_g N_VDD_Mp8@2706_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2705 N_OUT8_Mn8@2705_d N_OUT7_Mn8@2705_g N_VSS_Mn8@2705_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2704 N_OUT8_Mn8@2704_d N_OUT7_Mn8@2704_g N_VSS_Mn8@2704_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2705 N_OUT8_Mp8@2705_d N_OUT7_Mp8@2705_g N_VDD_Mp8@2705_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2704 N_OUT8_Mp8@2704_d N_OUT7_Mp8@2704_g N_VDD_Mp8@2704_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2703 N_OUT8_Mn8@2703_d N_OUT7_Mn8@2703_g N_VSS_Mn8@2703_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2702 N_OUT8_Mn8@2702_d N_OUT7_Mn8@2702_g N_VSS_Mn8@2702_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2703 N_OUT8_Mp8@2703_d N_OUT7_Mp8@2703_g N_VDD_Mp8@2703_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2702 N_OUT8_Mp8@2702_d N_OUT7_Mp8@2702_g N_VDD_Mp8@2702_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2701 N_OUT8_Mn8@2701_d N_OUT7_Mn8@2701_g N_VSS_Mn8@2701_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2700 N_OUT8_Mn8@2700_d N_OUT7_Mn8@2700_g N_VSS_Mn8@2700_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2701 N_OUT8_Mp8@2701_d N_OUT7_Mp8@2701_g N_VDD_Mp8@2701_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2700 N_OUT8_Mp8@2700_d N_OUT7_Mp8@2700_g N_VDD_Mp8@2700_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2699 N_OUT8_Mn8@2699_d N_OUT7_Mn8@2699_g N_VSS_Mn8@2699_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2698 N_OUT8_Mn8@2698_d N_OUT7_Mn8@2698_g N_VSS_Mn8@2698_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2699 N_OUT8_Mp8@2699_d N_OUT7_Mp8@2699_g N_VDD_Mp8@2699_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2698 N_OUT8_Mp8@2698_d N_OUT7_Mp8@2698_g N_VDD_Mp8@2698_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2697 N_OUT8_Mn8@2697_d N_OUT7_Mn8@2697_g N_VSS_Mn8@2697_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2696 N_OUT8_Mn8@2696_d N_OUT7_Mn8@2696_g N_VSS_Mn8@2696_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2697 N_OUT8_Mp8@2697_d N_OUT7_Mp8@2697_g N_VDD_Mp8@2697_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2696 N_OUT8_Mp8@2696_d N_OUT7_Mp8@2696_g N_VDD_Mp8@2696_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2695 N_OUT8_Mn8@2695_d N_OUT7_Mn8@2695_g N_VSS_Mn8@2695_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2694 N_OUT8_Mn8@2694_d N_OUT7_Mn8@2694_g N_VSS_Mn8@2694_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2695 N_OUT8_Mp8@2695_d N_OUT7_Mp8@2695_g N_VDD_Mp8@2695_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2694 N_OUT8_Mp8@2694_d N_OUT7_Mp8@2694_g N_VDD_Mp8@2694_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2693 N_OUT8_Mn8@2693_d N_OUT7_Mn8@2693_g N_VSS_Mn8@2693_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2692 N_OUT8_Mn8@2692_d N_OUT7_Mn8@2692_g N_VSS_Mn8@2692_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2693 N_OUT8_Mp8@2693_d N_OUT7_Mp8@2693_g N_VDD_Mp8@2693_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2692 N_OUT8_Mp8@2692_d N_OUT7_Mp8@2692_g N_VDD_Mp8@2692_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2691 N_OUT8_Mn8@2691_d N_OUT7_Mn8@2691_g N_VSS_Mn8@2691_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2690 N_OUT8_Mn8@2690_d N_OUT7_Mn8@2690_g N_VSS_Mn8@2690_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2691 N_OUT8_Mp8@2691_d N_OUT7_Mp8@2691_g N_VDD_Mp8@2691_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2690 N_OUT8_Mp8@2690_d N_OUT7_Mp8@2690_g N_VDD_Mp8@2690_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2689 N_OUT8_Mn8@2689_d N_OUT7_Mn8@2689_g N_VSS_Mn8@2689_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2688 N_OUT8_Mn8@2688_d N_OUT7_Mn8@2688_g N_VSS_Mn8@2688_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2689 N_OUT8_Mp8@2689_d N_OUT7_Mp8@2689_g N_VDD_Mp8@2689_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2688 N_OUT8_Mp8@2688_d N_OUT7_Mp8@2688_g N_VDD_Mp8@2688_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2687 N_OUT8_Mn8@2687_d N_OUT7_Mn8@2687_g N_VSS_Mn8@2687_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2686 N_OUT8_Mn8@2686_d N_OUT7_Mn8@2686_g N_VSS_Mn8@2686_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2687 N_OUT8_Mp8@2687_d N_OUT7_Mp8@2687_g N_VDD_Mp8@2687_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2686 N_OUT8_Mp8@2686_d N_OUT7_Mp8@2686_g N_VDD_Mp8@2686_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2685 N_OUT8_Mn8@2685_d N_OUT7_Mn8@2685_g N_VSS_Mn8@2685_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2684 N_OUT8_Mn8@2684_d N_OUT7_Mn8@2684_g N_VSS_Mn8@2684_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2685 N_OUT8_Mp8@2685_d N_OUT7_Mp8@2685_g N_VDD_Mp8@2685_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2684 N_OUT8_Mp8@2684_d N_OUT7_Mp8@2684_g N_VDD_Mp8@2684_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2683 N_OUT8_Mn8@2683_d N_OUT7_Mn8@2683_g N_VSS_Mn8@2683_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2682 N_OUT8_Mn8@2682_d N_OUT7_Mn8@2682_g N_VSS_Mn8@2682_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2683 N_OUT8_Mp8@2683_d N_OUT7_Mp8@2683_g N_VDD_Mp8@2683_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2682 N_OUT8_Mp8@2682_d N_OUT7_Mp8@2682_g N_VDD_Mp8@2682_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2681 N_OUT8_Mn8@2681_d N_OUT7_Mn8@2681_g N_VSS_Mn8@2681_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2680 N_OUT8_Mn8@2680_d N_OUT7_Mn8@2680_g N_VSS_Mn8@2680_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2681 N_OUT8_Mp8@2681_d N_OUT7_Mp8@2681_g N_VDD_Mp8@2681_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2680 N_OUT8_Mp8@2680_d N_OUT7_Mp8@2680_g N_VDD_Mp8@2680_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2679 N_OUT8_Mn8@2679_d N_OUT7_Mn8@2679_g N_VSS_Mn8@2679_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2678 N_OUT8_Mn8@2678_d N_OUT7_Mn8@2678_g N_VSS_Mn8@2678_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2679 N_OUT8_Mp8@2679_d N_OUT7_Mp8@2679_g N_VDD_Mp8@2679_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2678 N_OUT8_Mp8@2678_d N_OUT7_Mp8@2678_g N_VDD_Mp8@2678_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2677 N_OUT8_Mn8@2677_d N_OUT7_Mn8@2677_g N_VSS_Mn8@2677_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2676 N_OUT8_Mn8@2676_d N_OUT7_Mn8@2676_g N_VSS_Mn8@2676_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2677 N_OUT8_Mp8@2677_d N_OUT7_Mp8@2677_g N_VDD_Mp8@2677_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2676 N_OUT8_Mp8@2676_d N_OUT7_Mp8@2676_g N_VDD_Mp8@2676_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2675 N_OUT8_Mn8@2675_d N_OUT7_Mn8@2675_g N_VSS_Mn8@2675_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2674 N_OUT8_Mn8@2674_d N_OUT7_Mn8@2674_g N_VSS_Mn8@2674_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2675 N_OUT8_Mp8@2675_d N_OUT7_Mp8@2675_g N_VDD_Mp8@2675_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2674 N_OUT8_Mp8@2674_d N_OUT7_Mp8@2674_g N_VDD_Mp8@2674_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2673 N_OUT8_Mn8@2673_d N_OUT7_Mn8@2673_g N_VSS_Mn8@2673_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2672 N_OUT8_Mn8@2672_d N_OUT7_Mn8@2672_g N_VSS_Mn8@2672_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2673 N_OUT8_Mp8@2673_d N_OUT7_Mp8@2673_g N_VDD_Mp8@2673_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2672 N_OUT8_Mp8@2672_d N_OUT7_Mp8@2672_g N_VDD_Mp8@2672_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2671 N_OUT8_Mn8@2671_d N_OUT7_Mn8@2671_g N_VSS_Mn8@2671_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2670 N_OUT8_Mn8@2670_d N_OUT7_Mn8@2670_g N_VSS_Mn8@2670_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2671 N_OUT8_Mp8@2671_d N_OUT7_Mp8@2671_g N_VDD_Mp8@2671_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2670 N_OUT8_Mp8@2670_d N_OUT7_Mp8@2670_g N_VDD_Mp8@2670_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2669 N_OUT8_Mn8@2669_d N_OUT7_Mn8@2669_g N_VSS_Mn8@2669_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2668 N_OUT8_Mn8@2668_d N_OUT7_Mn8@2668_g N_VSS_Mn8@2668_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2669 N_OUT8_Mp8@2669_d N_OUT7_Mp8@2669_g N_VDD_Mp8@2669_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2668 N_OUT8_Mp8@2668_d N_OUT7_Mp8@2668_g N_VDD_Mp8@2668_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2667 N_OUT8_Mn8@2667_d N_OUT7_Mn8@2667_g N_VSS_Mn8@2667_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2666 N_OUT8_Mn8@2666_d N_OUT7_Mn8@2666_g N_VSS_Mn8@2666_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2667 N_OUT8_Mp8@2667_d N_OUT7_Mp8@2667_g N_VDD_Mp8@2667_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2666 N_OUT8_Mp8@2666_d N_OUT7_Mp8@2666_g N_VDD_Mp8@2666_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2665 N_OUT8_Mn8@2665_d N_OUT7_Mn8@2665_g N_VSS_Mn8@2665_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2664 N_OUT8_Mn8@2664_d N_OUT7_Mn8@2664_g N_VSS_Mn8@2664_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2665 N_OUT8_Mp8@2665_d N_OUT7_Mp8@2665_g N_VDD_Mp8@2665_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2664 N_OUT8_Mp8@2664_d N_OUT7_Mp8@2664_g N_VDD_Mp8@2664_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2663 N_OUT8_Mn8@2663_d N_OUT7_Mn8@2663_g N_VSS_Mn8@2663_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2662 N_OUT8_Mn8@2662_d N_OUT7_Mn8@2662_g N_VSS_Mn8@2662_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2663 N_OUT8_Mp8@2663_d N_OUT7_Mp8@2663_g N_VDD_Mp8@2663_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2662 N_OUT8_Mp8@2662_d N_OUT7_Mp8@2662_g N_VDD_Mp8@2662_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2661 N_OUT8_Mn8@2661_d N_OUT7_Mn8@2661_g N_VSS_Mn8@2661_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2660 N_OUT8_Mn8@2660_d N_OUT7_Mn8@2660_g N_VSS_Mn8@2660_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2661 N_OUT8_Mp8@2661_d N_OUT7_Mp8@2661_g N_VDD_Mp8@2661_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2660 N_OUT8_Mp8@2660_d N_OUT7_Mp8@2660_g N_VDD_Mp8@2660_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2659 N_OUT8_Mn8@2659_d N_OUT7_Mn8@2659_g N_VSS_Mn8@2659_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2658 N_OUT8_Mn8@2658_d N_OUT7_Mn8@2658_g N_VSS_Mn8@2658_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2659 N_OUT8_Mp8@2659_d N_OUT7_Mp8@2659_g N_VDD_Mp8@2659_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2658 N_OUT8_Mp8@2658_d N_OUT7_Mp8@2658_g N_VDD_Mp8@2658_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2657 N_OUT8_Mn8@2657_d N_OUT7_Mn8@2657_g N_VSS_Mn8@2657_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2656 N_OUT8_Mn8@2656_d N_OUT7_Mn8@2656_g N_VSS_Mn8@2656_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2657 N_OUT8_Mp8@2657_d N_OUT7_Mp8@2657_g N_VDD_Mp8@2657_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2656 N_OUT8_Mp8@2656_d N_OUT7_Mp8@2656_g N_VDD_Mp8@2656_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2655 N_OUT8_Mn8@2655_d N_OUT7_Mn8@2655_g N_VSS_Mn8@2655_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2654 N_OUT8_Mn8@2654_d N_OUT7_Mn8@2654_g N_VSS_Mn8@2654_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2655 N_OUT8_Mp8@2655_d N_OUT7_Mp8@2655_g N_VDD_Mp8@2655_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2654 N_OUT8_Mp8@2654_d N_OUT7_Mp8@2654_g N_VDD_Mp8@2654_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2653 N_OUT8_Mn8@2653_d N_OUT7_Mn8@2653_g N_VSS_Mn8@2653_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2652 N_OUT8_Mn8@2652_d N_OUT7_Mn8@2652_g N_VSS_Mn8@2652_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2653 N_OUT8_Mp8@2653_d N_OUT7_Mp8@2653_g N_VDD_Mp8@2653_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2652 N_OUT8_Mp8@2652_d N_OUT7_Mp8@2652_g N_VDD_Mp8@2652_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2651 N_OUT8_Mn8@2651_d N_OUT7_Mn8@2651_g N_VSS_Mn8@2651_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2650 N_OUT8_Mn8@2650_d N_OUT7_Mn8@2650_g N_VSS_Mn8@2650_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2651 N_OUT8_Mp8@2651_d N_OUT7_Mp8@2651_g N_VDD_Mp8@2651_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2650 N_OUT8_Mp8@2650_d N_OUT7_Mp8@2650_g N_VDD_Mp8@2650_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2649 N_OUT8_Mn8@2649_d N_OUT7_Mn8@2649_g N_VSS_Mn8@2649_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2648 N_OUT8_Mn8@2648_d N_OUT7_Mn8@2648_g N_VSS_Mn8@2648_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2649 N_OUT8_Mp8@2649_d N_OUT7_Mp8@2649_g N_VDD_Mp8@2649_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2648 N_OUT8_Mp8@2648_d N_OUT7_Mp8@2648_g N_VDD_Mp8@2648_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2647 N_OUT8_Mn8@2647_d N_OUT7_Mn8@2647_g N_VSS_Mn8@2647_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2646 N_OUT8_Mn8@2646_d N_OUT7_Mn8@2646_g N_VSS_Mn8@2646_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2647 N_OUT8_Mp8@2647_d N_OUT7_Mp8@2647_g N_VDD_Mp8@2647_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2646 N_OUT8_Mp8@2646_d N_OUT7_Mp8@2646_g N_VDD_Mp8@2646_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2645 N_OUT8_Mn8@2645_d N_OUT7_Mn8@2645_g N_VSS_Mn8@2645_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2644 N_OUT8_Mn8@2644_d N_OUT7_Mn8@2644_g N_VSS_Mn8@2644_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2645 N_OUT8_Mp8@2645_d N_OUT7_Mp8@2645_g N_VDD_Mp8@2645_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2644 N_OUT8_Mp8@2644_d N_OUT7_Mp8@2644_g N_VDD_Mp8@2644_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2643 N_OUT8_Mn8@2643_d N_OUT7_Mn8@2643_g N_VSS_Mn8@2643_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2642 N_OUT8_Mn8@2642_d N_OUT7_Mn8@2642_g N_VSS_Mn8@2642_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2643 N_OUT8_Mp8@2643_d N_OUT7_Mp8@2643_g N_VDD_Mp8@2643_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2642 N_OUT8_Mp8@2642_d N_OUT7_Mp8@2642_g N_VDD_Mp8@2642_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2641 N_OUT8_Mn8@2641_d N_OUT7_Mn8@2641_g N_VSS_Mn8@2641_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2640 N_OUT8_Mn8@2640_d N_OUT7_Mn8@2640_g N_VSS_Mn8@2640_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2641 N_OUT8_Mp8@2641_d N_OUT7_Mp8@2641_g N_VDD_Mp8@2641_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2640 N_OUT8_Mp8@2640_d N_OUT7_Mp8@2640_g N_VDD_Mp8@2640_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2639 N_OUT8_Mn8@2639_d N_OUT7_Mn8@2639_g N_VSS_Mn8@2639_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2638 N_OUT8_Mn8@2638_d N_OUT7_Mn8@2638_g N_VSS_Mn8@2638_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2639 N_OUT8_Mp8@2639_d N_OUT7_Mp8@2639_g N_VDD_Mp8@2639_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2638 N_OUT8_Mp8@2638_d N_OUT7_Mp8@2638_g N_VDD_Mp8@2638_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2637 N_OUT8_Mn8@2637_d N_OUT7_Mn8@2637_g N_VSS_Mn8@2637_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2636 N_OUT8_Mn8@2636_d N_OUT7_Mn8@2636_g N_VSS_Mn8@2636_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2637 N_OUT8_Mp8@2637_d N_OUT7_Mp8@2637_g N_VDD_Mp8@2637_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2636 N_OUT8_Mp8@2636_d N_OUT7_Mp8@2636_g N_VDD_Mp8@2636_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2635 N_OUT8_Mn8@2635_d N_OUT7_Mn8@2635_g N_VSS_Mn8@2635_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2634 N_OUT8_Mn8@2634_d N_OUT7_Mn8@2634_g N_VSS_Mn8@2634_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2635 N_OUT8_Mp8@2635_d N_OUT7_Mp8@2635_g N_VDD_Mp8@2635_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2634 N_OUT8_Mp8@2634_d N_OUT7_Mp8@2634_g N_VDD_Mp8@2634_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2633 N_OUT8_Mn8@2633_d N_OUT7_Mn8@2633_g N_VSS_Mn8@2633_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2632 N_OUT8_Mn8@2632_d N_OUT7_Mn8@2632_g N_VSS_Mn8@2632_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2633 N_OUT8_Mp8@2633_d N_OUT7_Mp8@2633_g N_VDD_Mp8@2633_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2632 N_OUT8_Mp8@2632_d N_OUT7_Mp8@2632_g N_VDD_Mp8@2632_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2631 N_OUT8_Mn8@2631_d N_OUT7_Mn8@2631_g N_VSS_Mn8@2631_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2630 N_OUT8_Mn8@2630_d N_OUT7_Mn8@2630_g N_VSS_Mn8@2630_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2631 N_OUT8_Mp8@2631_d N_OUT7_Mp8@2631_g N_VDD_Mp8@2631_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2630 N_OUT8_Mp8@2630_d N_OUT7_Mp8@2630_g N_VDD_Mp8@2630_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2629 N_OUT8_Mn8@2629_d N_OUT7_Mn8@2629_g N_VSS_Mn8@2629_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2628 N_OUT8_Mn8@2628_d N_OUT7_Mn8@2628_g N_VSS_Mn8@2628_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2629 N_OUT8_Mp8@2629_d N_OUT7_Mp8@2629_g N_VDD_Mp8@2629_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2628 N_OUT8_Mp8@2628_d N_OUT7_Mp8@2628_g N_VDD_Mp8@2628_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2627 N_OUT8_Mn8@2627_d N_OUT7_Mn8@2627_g N_VSS_Mn8@2627_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2626 N_OUT8_Mn8@2626_d N_OUT7_Mn8@2626_g N_VSS_Mn8@2626_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2627 N_OUT8_Mp8@2627_d N_OUT7_Mp8@2627_g N_VDD_Mp8@2627_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2626 N_OUT8_Mp8@2626_d N_OUT7_Mp8@2626_g N_VDD_Mp8@2626_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2625 N_OUT8_Mn8@2625_d N_OUT7_Mn8@2625_g N_VSS_Mn8@2625_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2624 N_OUT8_Mn8@2624_d N_OUT7_Mn8@2624_g N_VSS_Mn8@2624_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2625 N_OUT8_Mp8@2625_d N_OUT7_Mp8@2625_g N_VDD_Mp8@2625_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2624 N_OUT8_Mp8@2624_d N_OUT7_Mp8@2624_g N_VDD_Mp8@2624_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2623 N_OUT8_Mn8@2623_d N_OUT7_Mn8@2623_g N_VSS_Mn8@2623_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2622 N_OUT8_Mn8@2622_d N_OUT7_Mn8@2622_g N_VSS_Mn8@2622_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2623 N_OUT8_Mp8@2623_d N_OUT7_Mp8@2623_g N_VDD_Mp8@2623_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2622 N_OUT8_Mp8@2622_d N_OUT7_Mp8@2622_g N_VDD_Mp8@2622_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2621 N_OUT8_Mn8@2621_d N_OUT7_Mn8@2621_g N_VSS_Mn8@2621_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2620 N_OUT8_Mn8@2620_d N_OUT7_Mn8@2620_g N_VSS_Mn8@2620_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2621 N_OUT8_Mp8@2621_d N_OUT7_Mp8@2621_g N_VDD_Mp8@2621_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2620 N_OUT8_Mp8@2620_d N_OUT7_Mp8@2620_g N_VDD_Mp8@2620_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2619 N_OUT8_Mn8@2619_d N_OUT7_Mn8@2619_g N_VSS_Mn8@2619_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2618 N_OUT8_Mn8@2618_d N_OUT7_Mn8@2618_g N_VSS_Mn8@2618_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2619 N_OUT8_Mp8@2619_d N_OUT7_Mp8@2619_g N_VDD_Mp8@2619_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2618 N_OUT8_Mp8@2618_d N_OUT7_Mp8@2618_g N_VDD_Mp8@2618_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2617 N_OUT8_Mn8@2617_d N_OUT7_Mn8@2617_g N_VSS_Mn8@2617_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2616 N_OUT8_Mn8@2616_d N_OUT7_Mn8@2616_g N_VSS_Mn8@2616_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2617 N_OUT8_Mp8@2617_d N_OUT7_Mp8@2617_g N_VDD_Mp8@2617_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2616 N_OUT8_Mp8@2616_d N_OUT7_Mp8@2616_g N_VDD_Mp8@2616_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2615 N_OUT8_Mn8@2615_d N_OUT7_Mn8@2615_g N_VSS_Mn8@2615_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2614 N_OUT8_Mn8@2614_d N_OUT7_Mn8@2614_g N_VSS_Mn8@2614_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2615 N_OUT8_Mp8@2615_d N_OUT7_Mp8@2615_g N_VDD_Mp8@2615_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2614 N_OUT8_Mp8@2614_d N_OUT7_Mp8@2614_g N_VDD_Mp8@2614_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2613 N_OUT8_Mn8@2613_d N_OUT7_Mn8@2613_g N_VSS_Mn8@2613_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2612 N_OUT8_Mn8@2612_d N_OUT7_Mn8@2612_g N_VSS_Mn8@2612_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2613 N_OUT8_Mp8@2613_d N_OUT7_Mp8@2613_g N_VDD_Mp8@2613_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2612 N_OUT8_Mp8@2612_d N_OUT7_Mp8@2612_g N_VDD_Mp8@2612_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2611 N_OUT8_Mn8@2611_d N_OUT7_Mn8@2611_g N_VSS_Mn8@2611_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2610 N_OUT8_Mn8@2610_d N_OUT7_Mn8@2610_g N_VSS_Mn8@2610_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2611 N_OUT8_Mp8@2611_d N_OUT7_Mp8@2611_g N_VDD_Mp8@2611_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2610 N_OUT8_Mp8@2610_d N_OUT7_Mp8@2610_g N_VDD_Mp8@2610_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2609 N_OUT8_Mn8@2609_d N_OUT7_Mn8@2609_g N_VSS_Mn8@2609_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2608 N_OUT8_Mn8@2608_d N_OUT7_Mn8@2608_g N_VSS_Mn8@2608_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2609 N_OUT8_Mp8@2609_d N_OUT7_Mp8@2609_g N_VDD_Mp8@2609_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2608 N_OUT8_Mp8@2608_d N_OUT7_Mp8@2608_g N_VDD_Mp8@2608_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2607 N_OUT8_Mn8@2607_d N_OUT7_Mn8@2607_g N_VSS_Mn8@2607_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2606 N_OUT8_Mn8@2606_d N_OUT7_Mn8@2606_g N_VSS_Mn8@2606_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2607 N_OUT8_Mp8@2607_d N_OUT7_Mp8@2607_g N_VDD_Mp8@2607_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2606 N_OUT8_Mp8@2606_d N_OUT7_Mp8@2606_g N_VDD_Mp8@2606_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2605 N_OUT8_Mn8@2605_d N_OUT7_Mn8@2605_g N_VSS_Mn8@2605_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2604 N_OUT8_Mn8@2604_d N_OUT7_Mn8@2604_g N_VSS_Mn8@2604_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2605 N_OUT8_Mp8@2605_d N_OUT7_Mp8@2605_g N_VDD_Mp8@2605_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2604 N_OUT8_Mp8@2604_d N_OUT7_Mp8@2604_g N_VDD_Mp8@2604_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2603 N_OUT8_Mn8@2603_d N_OUT7_Mn8@2603_g N_VSS_Mn8@2603_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2602 N_OUT8_Mn8@2602_d N_OUT7_Mn8@2602_g N_VSS_Mn8@2602_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2603 N_OUT8_Mp8@2603_d N_OUT7_Mp8@2603_g N_VDD_Mp8@2603_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2602 N_OUT8_Mp8@2602_d N_OUT7_Mp8@2602_g N_VDD_Mp8@2602_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2601 N_OUT8_Mn8@2601_d N_OUT7_Mn8@2601_g N_VSS_Mn8@2601_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2600 N_OUT8_Mn8@2600_d N_OUT7_Mn8@2600_g N_VSS_Mn8@2600_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2601 N_OUT8_Mp8@2601_d N_OUT7_Mp8@2601_g N_VDD_Mp8@2601_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2600 N_OUT8_Mp8@2600_d N_OUT7_Mp8@2600_g N_VDD_Mp8@2600_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2599 N_OUT8_Mn8@2599_d N_OUT7_Mn8@2599_g N_VSS_Mn8@2599_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2598 N_OUT8_Mn8@2598_d N_OUT7_Mn8@2598_g N_VSS_Mn8@2598_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2599 N_OUT8_Mp8@2599_d N_OUT7_Mp8@2599_g N_VDD_Mp8@2599_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2598 N_OUT8_Mp8@2598_d N_OUT7_Mp8@2598_g N_VDD_Mp8@2598_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2597 N_OUT8_Mn8@2597_d N_OUT7_Mn8@2597_g N_VSS_Mn8@2597_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2596 N_OUT8_Mn8@2596_d N_OUT7_Mn8@2596_g N_VSS_Mn8@2596_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2597 N_OUT8_Mp8@2597_d N_OUT7_Mp8@2597_g N_VDD_Mp8@2597_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2596 N_OUT8_Mp8@2596_d N_OUT7_Mp8@2596_g N_VDD_Mp8@2596_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2595 N_OUT8_Mn8@2595_d N_OUT7_Mn8@2595_g N_VSS_Mn8@2595_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2594 N_OUT8_Mn8@2594_d N_OUT7_Mn8@2594_g N_VSS_Mn8@2594_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2595 N_OUT8_Mp8@2595_d N_OUT7_Mp8@2595_g N_VDD_Mp8@2595_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2594 N_OUT8_Mp8@2594_d N_OUT7_Mp8@2594_g N_VDD_Mp8@2594_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2593 N_OUT8_Mn8@2593_d N_OUT7_Mn8@2593_g N_VSS_Mn8@2593_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2592 N_OUT8_Mn8@2592_d N_OUT7_Mn8@2592_g N_VSS_Mn8@2592_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2593 N_OUT8_Mp8@2593_d N_OUT7_Mp8@2593_g N_VDD_Mp8@2593_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2592 N_OUT8_Mp8@2592_d N_OUT7_Mp8@2592_g N_VDD_Mp8@2592_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2591 N_OUT8_Mn8@2591_d N_OUT7_Mn8@2591_g N_VSS_Mn8@2591_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2590 N_OUT8_Mn8@2590_d N_OUT7_Mn8@2590_g N_VSS_Mn8@2590_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2591 N_OUT8_Mp8@2591_d N_OUT7_Mp8@2591_g N_VDD_Mp8@2591_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2590 N_OUT8_Mp8@2590_d N_OUT7_Mp8@2590_g N_VDD_Mp8@2590_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2589 N_OUT8_Mn8@2589_d N_OUT7_Mn8@2589_g N_VSS_Mn8@2589_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2588 N_OUT8_Mn8@2588_d N_OUT7_Mn8@2588_g N_VSS_Mn8@2588_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2589 N_OUT8_Mp8@2589_d N_OUT7_Mp8@2589_g N_VDD_Mp8@2589_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2588 N_OUT8_Mp8@2588_d N_OUT7_Mp8@2588_g N_VDD_Mp8@2588_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2587 N_OUT8_Mn8@2587_d N_OUT7_Mn8@2587_g N_VSS_Mn8@2587_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2586 N_OUT8_Mn8@2586_d N_OUT7_Mn8@2586_g N_VSS_Mn8@2586_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2587 N_OUT8_Mp8@2587_d N_OUT7_Mp8@2587_g N_VDD_Mp8@2587_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2586 N_OUT8_Mp8@2586_d N_OUT7_Mp8@2586_g N_VDD_Mp8@2586_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2585 N_OUT8_Mn8@2585_d N_OUT7_Mn8@2585_g N_VSS_Mn8@2585_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2584 N_OUT8_Mn8@2584_d N_OUT7_Mn8@2584_g N_VSS_Mn8@2584_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2585 N_OUT8_Mp8@2585_d N_OUT7_Mp8@2585_g N_VDD_Mp8@2585_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2584 N_OUT8_Mp8@2584_d N_OUT7_Mp8@2584_g N_VDD_Mp8@2584_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2583 N_OUT8_Mn8@2583_d N_OUT7_Mn8@2583_g N_VSS_Mn8@2583_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2582 N_OUT8_Mn8@2582_d N_OUT7_Mn8@2582_g N_VSS_Mn8@2582_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2583 N_OUT8_Mp8@2583_d N_OUT7_Mp8@2583_g N_VDD_Mp8@2583_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2582 N_OUT8_Mp8@2582_d N_OUT7_Mp8@2582_g N_VDD_Mp8@2582_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2581 N_OUT8_Mn8@2581_d N_OUT7_Mn8@2581_g N_VSS_Mn8@2581_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2580 N_OUT8_Mn8@2580_d N_OUT7_Mn8@2580_g N_VSS_Mn8@2580_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2581 N_OUT8_Mp8@2581_d N_OUT7_Mp8@2581_g N_VDD_Mp8@2581_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2580 N_OUT8_Mp8@2580_d N_OUT7_Mp8@2580_g N_VDD_Mp8@2580_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2579 N_OUT8_Mn8@2579_d N_OUT7_Mn8@2579_g N_VSS_Mn8@2579_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2578 N_OUT8_Mn8@2578_d N_OUT7_Mn8@2578_g N_VSS_Mn8@2578_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2579 N_OUT8_Mp8@2579_d N_OUT7_Mp8@2579_g N_VDD_Mp8@2579_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2578 N_OUT8_Mp8@2578_d N_OUT7_Mp8@2578_g N_VDD_Mp8@2578_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2577 N_OUT8_Mn8@2577_d N_OUT7_Mn8@2577_g N_VSS_Mn8@2577_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2576 N_OUT8_Mn8@2576_d N_OUT7_Mn8@2576_g N_VSS_Mn8@2576_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2577 N_OUT8_Mp8@2577_d N_OUT7_Mp8@2577_g N_VDD_Mp8@2577_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2576 N_OUT8_Mp8@2576_d N_OUT7_Mp8@2576_g N_VDD_Mp8@2576_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2575 N_OUT8_Mn8@2575_d N_OUT7_Mn8@2575_g N_VSS_Mn8@2575_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2574 N_OUT8_Mn8@2574_d N_OUT7_Mn8@2574_g N_VSS_Mn8@2574_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2575 N_OUT8_Mp8@2575_d N_OUT7_Mp8@2575_g N_VDD_Mp8@2575_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2574 N_OUT8_Mp8@2574_d N_OUT7_Mp8@2574_g N_VDD_Mp8@2574_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2573 N_OUT8_Mn8@2573_d N_OUT7_Mn8@2573_g N_VSS_Mn8@2573_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2572 N_OUT8_Mn8@2572_d N_OUT7_Mn8@2572_g N_VSS_Mn8@2572_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2573 N_OUT8_Mp8@2573_d N_OUT7_Mp8@2573_g N_VDD_Mp8@2573_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2572 N_OUT8_Mp8@2572_d N_OUT7_Mp8@2572_g N_VDD_Mp8@2572_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2571 N_OUT8_Mn8@2571_d N_OUT7_Mn8@2571_g N_VSS_Mn8@2571_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2570 N_OUT8_Mn8@2570_d N_OUT7_Mn8@2570_g N_VSS_Mn8@2570_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2571 N_OUT8_Mp8@2571_d N_OUT7_Mp8@2571_g N_VDD_Mp8@2571_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2570 N_OUT8_Mp8@2570_d N_OUT7_Mp8@2570_g N_VDD_Mp8@2570_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2569 N_OUT8_Mn8@2569_d N_OUT7_Mn8@2569_g N_VSS_Mn8@2569_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2568 N_OUT8_Mn8@2568_d N_OUT7_Mn8@2568_g N_VSS_Mn8@2568_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2569 N_OUT8_Mp8@2569_d N_OUT7_Mp8@2569_g N_VDD_Mp8@2569_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2568 N_OUT8_Mp8@2568_d N_OUT7_Mp8@2568_g N_VDD_Mp8@2568_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2567 N_OUT8_Mn8@2567_d N_OUT7_Mn8@2567_g N_VSS_Mn8@2567_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2566 N_OUT8_Mn8@2566_d N_OUT7_Mn8@2566_g N_VSS_Mn8@2566_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2567 N_OUT8_Mp8@2567_d N_OUT7_Mp8@2567_g N_VDD_Mp8@2567_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2566 N_OUT8_Mp8@2566_d N_OUT7_Mp8@2566_g N_VDD_Mp8@2566_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2565 N_OUT8_Mn8@2565_d N_OUT7_Mn8@2565_g N_VSS_Mn8@2565_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2564 N_OUT8_Mn8@2564_d N_OUT7_Mn8@2564_g N_VSS_Mn8@2564_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2565 N_OUT8_Mp8@2565_d N_OUT7_Mp8@2565_g N_VDD_Mp8@2565_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2564 N_OUT8_Mp8@2564_d N_OUT7_Mp8@2564_g N_VDD_Mp8@2564_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2563 N_OUT8_Mn8@2563_d N_OUT7_Mn8@2563_g N_VSS_Mn8@2563_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2562 N_OUT8_Mn8@2562_d N_OUT7_Mn8@2562_g N_VSS_Mn8@2562_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2563 N_OUT8_Mp8@2563_d N_OUT7_Mp8@2563_g N_VDD_Mp8@2563_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2562 N_OUT8_Mp8@2562_d N_OUT7_Mp8@2562_g N_VDD_Mp8@2562_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2561 N_OUT8_Mn8@2561_d N_OUT7_Mn8@2561_g N_VSS_Mn8@2561_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2560 N_OUT8_Mn8@2560_d N_OUT7_Mn8@2560_g N_VSS_Mn8@2560_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2561 N_OUT8_Mp8@2561_d N_OUT7_Mp8@2561_g N_VDD_Mp8@2561_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2560 N_OUT8_Mp8@2560_d N_OUT7_Mp8@2560_g N_VDD_Mp8@2560_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2559 N_OUT8_Mn8@2559_d N_OUT7_Mn8@2559_g N_VSS_Mn8@2559_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2558 N_OUT8_Mn8@2558_d N_OUT7_Mn8@2558_g N_VSS_Mn8@2558_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2559 N_OUT8_Mp8@2559_d N_OUT7_Mp8@2559_g N_VDD_Mp8@2559_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2558 N_OUT8_Mp8@2558_d N_OUT7_Mp8@2558_g N_VDD_Mp8@2558_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2557 N_OUT8_Mn8@2557_d N_OUT7_Mn8@2557_g N_VSS_Mn8@2557_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2556 N_OUT8_Mn8@2556_d N_OUT7_Mn8@2556_g N_VSS_Mn8@2556_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2557 N_OUT8_Mp8@2557_d N_OUT7_Mp8@2557_g N_VDD_Mp8@2557_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2556 N_OUT8_Mp8@2556_d N_OUT7_Mp8@2556_g N_VDD_Mp8@2556_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2555 N_OUT8_Mn8@2555_d N_OUT7_Mn8@2555_g N_VSS_Mn8@2555_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2554 N_OUT8_Mn8@2554_d N_OUT7_Mn8@2554_g N_VSS_Mn8@2554_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2555 N_OUT8_Mp8@2555_d N_OUT7_Mp8@2555_g N_VDD_Mp8@2555_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2554 N_OUT8_Mp8@2554_d N_OUT7_Mp8@2554_g N_VDD_Mp8@2554_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2553 N_OUT8_Mn8@2553_d N_OUT7_Mn8@2553_g N_VSS_Mn8@2553_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2552 N_OUT8_Mn8@2552_d N_OUT7_Mn8@2552_g N_VSS_Mn8@2552_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2553 N_OUT8_Mp8@2553_d N_OUT7_Mp8@2553_g N_VDD_Mp8@2553_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2552 N_OUT8_Mp8@2552_d N_OUT7_Mp8@2552_g N_VDD_Mp8@2552_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2551 N_OUT8_Mn8@2551_d N_OUT7_Mn8@2551_g N_VSS_Mn8@2551_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2550 N_OUT8_Mn8@2550_d N_OUT7_Mn8@2550_g N_VSS_Mn8@2550_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2551 N_OUT8_Mp8@2551_d N_OUT7_Mp8@2551_g N_VDD_Mp8@2551_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2550 N_OUT8_Mp8@2550_d N_OUT7_Mp8@2550_g N_VDD_Mp8@2550_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2549 N_OUT8_Mn8@2549_d N_OUT7_Mn8@2549_g N_VSS_Mn8@2549_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2548 N_OUT8_Mn8@2548_d N_OUT7_Mn8@2548_g N_VSS_Mn8@2548_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2549 N_OUT8_Mp8@2549_d N_OUT7_Mp8@2549_g N_VDD_Mp8@2549_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2548 N_OUT8_Mp8@2548_d N_OUT7_Mp8@2548_g N_VDD_Mp8@2548_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2547 N_OUT8_Mn8@2547_d N_OUT7_Mn8@2547_g N_VSS_Mn8@2547_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2546 N_OUT8_Mn8@2546_d N_OUT7_Mn8@2546_g N_VSS_Mn8@2546_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2547 N_OUT8_Mp8@2547_d N_OUT7_Mp8@2547_g N_VDD_Mp8@2547_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2546 N_OUT8_Mp8@2546_d N_OUT7_Mp8@2546_g N_VDD_Mp8@2546_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2545 N_OUT8_Mn8@2545_d N_OUT7_Mn8@2545_g N_VSS_Mn8@2545_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2544 N_OUT8_Mn8@2544_d N_OUT7_Mn8@2544_g N_VSS_Mn8@2544_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2545 N_OUT8_Mp8@2545_d N_OUT7_Mp8@2545_g N_VDD_Mp8@2545_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2544 N_OUT8_Mp8@2544_d N_OUT7_Mp8@2544_g N_VDD_Mp8@2544_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2543 N_OUT8_Mn8@2543_d N_OUT7_Mn8@2543_g N_VSS_Mn8@2543_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2542 N_OUT8_Mn8@2542_d N_OUT7_Mn8@2542_g N_VSS_Mn8@2542_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2543 N_OUT8_Mp8@2543_d N_OUT7_Mp8@2543_g N_VDD_Mp8@2543_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2542 N_OUT8_Mp8@2542_d N_OUT7_Mp8@2542_g N_VDD_Mp8@2542_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2541 N_OUT8_Mn8@2541_d N_OUT7_Mn8@2541_g N_VSS_Mn8@2541_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2540 N_OUT8_Mn8@2540_d N_OUT7_Mn8@2540_g N_VSS_Mn8@2540_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2541 N_OUT8_Mp8@2541_d N_OUT7_Mp8@2541_g N_VDD_Mp8@2541_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2540 N_OUT8_Mp8@2540_d N_OUT7_Mp8@2540_g N_VDD_Mp8@2540_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2539 N_OUT8_Mn8@2539_d N_OUT7_Mn8@2539_g N_VSS_Mn8@2539_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2538 N_OUT8_Mn8@2538_d N_OUT7_Mn8@2538_g N_VSS_Mn8@2538_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2539 N_OUT8_Mp8@2539_d N_OUT7_Mp8@2539_g N_VDD_Mp8@2539_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2538 N_OUT8_Mp8@2538_d N_OUT7_Mp8@2538_g N_VDD_Mp8@2538_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2537 N_OUT8_Mn8@2537_d N_OUT7_Mn8@2537_g N_VSS_Mn8@2537_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2536 N_OUT8_Mn8@2536_d N_OUT7_Mn8@2536_g N_VSS_Mn8@2536_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2537 N_OUT8_Mp8@2537_d N_OUT7_Mp8@2537_g N_VDD_Mp8@2537_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2536 N_OUT8_Mp8@2536_d N_OUT7_Mp8@2536_g N_VDD_Mp8@2536_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2535 N_OUT8_Mn8@2535_d N_OUT7_Mn8@2535_g N_VSS_Mn8@2535_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2534 N_OUT8_Mn8@2534_d N_OUT7_Mn8@2534_g N_VSS_Mn8@2534_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2535 N_OUT8_Mp8@2535_d N_OUT7_Mp8@2535_g N_VDD_Mp8@2535_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2534 N_OUT8_Mp8@2534_d N_OUT7_Mp8@2534_g N_VDD_Mp8@2534_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2533 N_OUT8_Mn8@2533_d N_OUT7_Mn8@2533_g N_VSS_Mn8@2533_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2532 N_OUT8_Mn8@2532_d N_OUT7_Mn8@2532_g N_VSS_Mn8@2532_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2533 N_OUT8_Mp8@2533_d N_OUT7_Mp8@2533_g N_VDD_Mp8@2533_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2532 N_OUT8_Mp8@2532_d N_OUT7_Mp8@2532_g N_VDD_Mp8@2532_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2531 N_OUT8_Mn8@2531_d N_OUT7_Mn8@2531_g N_VSS_Mn8@2531_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2530 N_OUT8_Mn8@2530_d N_OUT7_Mn8@2530_g N_VSS_Mn8@2530_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2531 N_OUT8_Mp8@2531_d N_OUT7_Mp8@2531_g N_VDD_Mp8@2531_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2530 N_OUT8_Mp8@2530_d N_OUT7_Mp8@2530_g N_VDD_Mp8@2530_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2529 N_OUT8_Mn8@2529_d N_OUT7_Mn8@2529_g N_VSS_Mn8@2529_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2528 N_OUT8_Mn8@2528_d N_OUT7_Mn8@2528_g N_VSS_Mn8@2528_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2529 N_OUT8_Mp8@2529_d N_OUT7_Mp8@2529_g N_VDD_Mp8@2529_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2528 N_OUT8_Mp8@2528_d N_OUT7_Mp8@2528_g N_VDD_Mp8@2528_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2527 N_OUT8_Mn8@2527_d N_OUT7_Mn8@2527_g N_VSS_Mn8@2527_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2526 N_OUT8_Mn8@2526_d N_OUT7_Mn8@2526_g N_VSS_Mn8@2526_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2527 N_OUT8_Mp8@2527_d N_OUT7_Mp8@2527_g N_VDD_Mp8@2527_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2526 N_OUT8_Mp8@2526_d N_OUT7_Mp8@2526_g N_VDD_Mp8@2526_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2525 N_OUT8_Mn8@2525_d N_OUT7_Mn8@2525_g N_VSS_Mn8@2525_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2524 N_OUT8_Mn8@2524_d N_OUT7_Mn8@2524_g N_VSS_Mn8@2524_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2525 N_OUT8_Mp8@2525_d N_OUT7_Mp8@2525_g N_VDD_Mp8@2525_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2524 N_OUT8_Mp8@2524_d N_OUT7_Mp8@2524_g N_VDD_Mp8@2524_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2523 N_OUT8_Mn8@2523_d N_OUT7_Mn8@2523_g N_VSS_Mn8@2523_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2522 N_OUT8_Mn8@2522_d N_OUT7_Mn8@2522_g N_VSS_Mn8@2522_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2523 N_OUT8_Mp8@2523_d N_OUT7_Mp8@2523_g N_VDD_Mp8@2523_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2522 N_OUT8_Mp8@2522_d N_OUT7_Mp8@2522_g N_VDD_Mp8@2522_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2521 N_OUT8_Mn8@2521_d N_OUT7_Mn8@2521_g N_VSS_Mn8@2521_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2520 N_OUT8_Mn8@2520_d N_OUT7_Mn8@2520_g N_VSS_Mn8@2520_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2521 N_OUT8_Mp8@2521_d N_OUT7_Mp8@2521_g N_VDD_Mp8@2521_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2520 N_OUT8_Mp8@2520_d N_OUT7_Mp8@2520_g N_VDD_Mp8@2520_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2519 N_OUT8_Mn8@2519_d N_OUT7_Mn8@2519_g N_VSS_Mn8@2519_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2518 N_OUT8_Mn8@2518_d N_OUT7_Mn8@2518_g N_VSS_Mn8@2518_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2519 N_OUT8_Mp8@2519_d N_OUT7_Mp8@2519_g N_VDD_Mp8@2519_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2518 N_OUT8_Mp8@2518_d N_OUT7_Mp8@2518_g N_VDD_Mp8@2518_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2517 N_OUT8_Mn8@2517_d N_OUT7_Mn8@2517_g N_VSS_Mn8@2517_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2516 N_OUT8_Mn8@2516_d N_OUT7_Mn8@2516_g N_VSS_Mn8@2516_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2517 N_OUT8_Mp8@2517_d N_OUT7_Mp8@2517_g N_VDD_Mp8@2517_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2516 N_OUT8_Mp8@2516_d N_OUT7_Mp8@2516_g N_VDD_Mp8@2516_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2515 N_OUT8_Mn8@2515_d N_OUT7_Mn8@2515_g N_VSS_Mn8@2515_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2514 N_OUT8_Mn8@2514_d N_OUT7_Mn8@2514_g N_VSS_Mn8@2514_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2515 N_OUT8_Mp8@2515_d N_OUT7_Mp8@2515_g N_VDD_Mp8@2515_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2514 N_OUT8_Mp8@2514_d N_OUT7_Mp8@2514_g N_VDD_Mp8@2514_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2513 N_OUT8_Mn8@2513_d N_OUT7_Mn8@2513_g N_VSS_Mn8@2513_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2512 N_OUT8_Mn8@2512_d N_OUT7_Mn8@2512_g N_VSS_Mn8@2512_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2513 N_OUT8_Mp8@2513_d N_OUT7_Mp8@2513_g N_VDD_Mp8@2513_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2512 N_OUT8_Mp8@2512_d N_OUT7_Mp8@2512_g N_VDD_Mp8@2512_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2511 N_OUT8_Mn8@2511_d N_OUT7_Mn8@2511_g N_VSS_Mn8@2511_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2510 N_OUT8_Mn8@2510_d N_OUT7_Mn8@2510_g N_VSS_Mn8@2510_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2511 N_OUT8_Mp8@2511_d N_OUT7_Mp8@2511_g N_VDD_Mp8@2511_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2510 N_OUT8_Mp8@2510_d N_OUT7_Mp8@2510_g N_VDD_Mp8@2510_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2509 N_OUT8_Mn8@2509_d N_OUT7_Mn8@2509_g N_VSS_Mn8@2509_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2508 N_OUT8_Mn8@2508_d N_OUT7_Mn8@2508_g N_VSS_Mn8@2508_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2509 N_OUT8_Mp8@2509_d N_OUT7_Mp8@2509_g N_VDD_Mp8@2509_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2508 N_OUT8_Mp8@2508_d N_OUT7_Mp8@2508_g N_VDD_Mp8@2508_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2507 N_OUT8_Mn8@2507_d N_OUT7_Mn8@2507_g N_VSS_Mn8@2507_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2506 N_OUT8_Mn8@2506_d N_OUT7_Mn8@2506_g N_VSS_Mn8@2506_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2507 N_OUT8_Mp8@2507_d N_OUT7_Mp8@2507_g N_VDD_Mp8@2507_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2506 N_OUT8_Mp8@2506_d N_OUT7_Mp8@2506_g N_VDD_Mp8@2506_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2505 N_OUT8_Mn8@2505_d N_OUT7_Mn8@2505_g N_VSS_Mn8@2505_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2504 N_OUT8_Mn8@2504_d N_OUT7_Mn8@2504_g N_VSS_Mn8@2504_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2505 N_OUT8_Mp8@2505_d N_OUT7_Mp8@2505_g N_VDD_Mp8@2505_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2504 N_OUT8_Mp8@2504_d N_OUT7_Mp8@2504_g N_VDD_Mp8@2504_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2503 N_OUT8_Mn8@2503_d N_OUT7_Mn8@2503_g N_VSS_Mn8@2503_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2502 N_OUT8_Mn8@2502_d N_OUT7_Mn8@2502_g N_VSS_Mn8@2502_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2503 N_OUT8_Mp8@2503_d N_OUT7_Mp8@2503_g N_VDD_Mp8@2503_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2502 N_OUT8_Mp8@2502_d N_OUT7_Mp8@2502_g N_VDD_Mp8@2502_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2501 N_OUT8_Mn8@2501_d N_OUT7_Mn8@2501_g N_VSS_Mn8@2501_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2500 N_OUT8_Mn8@2500_d N_OUT7_Mn8@2500_g N_VSS_Mn8@2500_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2501 N_OUT8_Mp8@2501_d N_OUT7_Mp8@2501_g N_VDD_Mp8@2501_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2500 N_OUT8_Mp8@2500_d N_OUT7_Mp8@2500_g N_VDD_Mp8@2500_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2499 N_OUT8_Mn8@2499_d N_OUT7_Mn8@2499_g N_VSS_Mn8@2499_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2498 N_OUT8_Mn8@2498_d N_OUT7_Mn8@2498_g N_VSS_Mn8@2498_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2499 N_OUT8_Mp8@2499_d N_OUT7_Mp8@2499_g N_VDD_Mp8@2499_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2498 N_OUT8_Mp8@2498_d N_OUT7_Mp8@2498_g N_VDD_Mp8@2498_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2497 N_OUT8_Mn8@2497_d N_OUT7_Mn8@2497_g N_VSS_Mn8@2497_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2496 N_OUT8_Mn8@2496_d N_OUT7_Mn8@2496_g N_VSS_Mn8@2496_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2497 N_OUT8_Mp8@2497_d N_OUT7_Mp8@2497_g N_VDD_Mp8@2497_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2496 N_OUT8_Mp8@2496_d N_OUT7_Mp8@2496_g N_VDD_Mp8@2496_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2495 N_OUT8_Mn8@2495_d N_OUT7_Mn8@2495_g N_VSS_Mn8@2495_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2494 N_OUT8_Mn8@2494_d N_OUT7_Mn8@2494_g N_VSS_Mn8@2494_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2495 N_OUT8_Mp8@2495_d N_OUT7_Mp8@2495_g N_VDD_Mp8@2495_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2494 N_OUT8_Mp8@2494_d N_OUT7_Mp8@2494_g N_VDD_Mp8@2494_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2493 N_OUT8_Mn8@2493_d N_OUT7_Mn8@2493_g N_VSS_Mn8@2493_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2492 N_OUT8_Mn8@2492_d N_OUT7_Mn8@2492_g N_VSS_Mn8@2492_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2493 N_OUT8_Mp8@2493_d N_OUT7_Mp8@2493_g N_VDD_Mp8@2493_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2492 N_OUT8_Mp8@2492_d N_OUT7_Mp8@2492_g N_VDD_Mp8@2492_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2491 N_OUT8_Mn8@2491_d N_OUT7_Mn8@2491_g N_VSS_Mn8@2491_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2490 N_OUT8_Mn8@2490_d N_OUT7_Mn8@2490_g N_VSS_Mn8@2490_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2491 N_OUT8_Mp8@2491_d N_OUT7_Mp8@2491_g N_VDD_Mp8@2491_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2490 N_OUT8_Mp8@2490_d N_OUT7_Mp8@2490_g N_VDD_Mp8@2490_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2489 N_OUT8_Mn8@2489_d N_OUT7_Mn8@2489_g N_VSS_Mn8@2489_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2488 N_OUT8_Mn8@2488_d N_OUT7_Mn8@2488_g N_VSS_Mn8@2488_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2489 N_OUT8_Mp8@2489_d N_OUT7_Mp8@2489_g N_VDD_Mp8@2489_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2488 N_OUT8_Mp8@2488_d N_OUT7_Mp8@2488_g N_VDD_Mp8@2488_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2487 N_OUT8_Mn8@2487_d N_OUT7_Mn8@2487_g N_VSS_Mn8@2487_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2486 N_OUT8_Mn8@2486_d N_OUT7_Mn8@2486_g N_VSS_Mn8@2486_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2487 N_OUT8_Mp8@2487_d N_OUT7_Mp8@2487_g N_VDD_Mp8@2487_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2486 N_OUT8_Mp8@2486_d N_OUT7_Mp8@2486_g N_VDD_Mp8@2486_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2485 N_OUT8_Mn8@2485_d N_OUT7_Mn8@2485_g N_VSS_Mn8@2485_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2484 N_OUT8_Mn8@2484_d N_OUT7_Mn8@2484_g N_VSS_Mn8@2484_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2485 N_OUT8_Mp8@2485_d N_OUT7_Mp8@2485_g N_VDD_Mp8@2485_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2484 N_OUT8_Mp8@2484_d N_OUT7_Mp8@2484_g N_VDD_Mp8@2484_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2483 N_OUT8_Mn8@2483_d N_OUT7_Mn8@2483_g N_VSS_Mn8@2483_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2482 N_OUT8_Mn8@2482_d N_OUT7_Mn8@2482_g N_VSS_Mn8@2482_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2483 N_OUT8_Mp8@2483_d N_OUT7_Mp8@2483_g N_VDD_Mp8@2483_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2482 N_OUT8_Mp8@2482_d N_OUT7_Mp8@2482_g N_VDD_Mp8@2482_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2481 N_OUT8_Mn8@2481_d N_OUT7_Mn8@2481_g N_VSS_Mn8@2481_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2480 N_OUT8_Mn8@2480_d N_OUT7_Mn8@2480_g N_VSS_Mn8@2480_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2481 N_OUT8_Mp8@2481_d N_OUT7_Mp8@2481_g N_VDD_Mp8@2481_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2480 N_OUT8_Mp8@2480_d N_OUT7_Mp8@2480_g N_VDD_Mp8@2480_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2479 N_OUT8_Mn8@2479_d N_OUT7_Mn8@2479_g N_VSS_Mn8@2479_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2478 N_OUT8_Mn8@2478_d N_OUT7_Mn8@2478_g N_VSS_Mn8@2478_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2479 N_OUT8_Mp8@2479_d N_OUT7_Mp8@2479_g N_VDD_Mp8@2479_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2478 N_OUT8_Mp8@2478_d N_OUT7_Mp8@2478_g N_VDD_Mp8@2478_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2477 N_OUT8_Mn8@2477_d N_OUT7_Mn8@2477_g N_VSS_Mn8@2477_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2476 N_OUT8_Mn8@2476_d N_OUT7_Mn8@2476_g N_VSS_Mn8@2476_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2477 N_OUT8_Mp8@2477_d N_OUT7_Mp8@2477_g N_VDD_Mp8@2477_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2476 N_OUT8_Mp8@2476_d N_OUT7_Mp8@2476_g N_VDD_Mp8@2476_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2475 N_OUT8_Mn8@2475_d N_OUT7_Mn8@2475_g N_VSS_Mn8@2475_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2474 N_OUT8_Mn8@2474_d N_OUT7_Mn8@2474_g N_VSS_Mn8@2474_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2475 N_OUT8_Mp8@2475_d N_OUT7_Mp8@2475_g N_VDD_Mp8@2475_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2474 N_OUT8_Mp8@2474_d N_OUT7_Mp8@2474_g N_VDD_Mp8@2474_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2473 N_OUT8_Mn8@2473_d N_OUT7_Mn8@2473_g N_VSS_Mn8@2473_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2472 N_OUT8_Mn8@2472_d N_OUT7_Mn8@2472_g N_VSS_Mn8@2472_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2473 N_OUT8_Mp8@2473_d N_OUT7_Mp8@2473_g N_VDD_Mp8@2473_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2472 N_OUT8_Mp8@2472_d N_OUT7_Mp8@2472_g N_VDD_Mp8@2472_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2471 N_OUT8_Mn8@2471_d N_OUT7_Mn8@2471_g N_VSS_Mn8@2471_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2470 N_OUT8_Mn8@2470_d N_OUT7_Mn8@2470_g N_VSS_Mn8@2470_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2471 N_OUT8_Mp8@2471_d N_OUT7_Mp8@2471_g N_VDD_Mp8@2471_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2470 N_OUT8_Mp8@2470_d N_OUT7_Mp8@2470_g N_VDD_Mp8@2470_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2469 N_OUT8_Mn8@2469_d N_OUT7_Mn8@2469_g N_VSS_Mn8@2469_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2468 N_OUT8_Mn8@2468_d N_OUT7_Mn8@2468_g N_VSS_Mn8@2468_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2469 N_OUT8_Mp8@2469_d N_OUT7_Mp8@2469_g N_VDD_Mp8@2469_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2468 N_OUT8_Mp8@2468_d N_OUT7_Mp8@2468_g N_VDD_Mp8@2468_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2467 N_OUT8_Mn8@2467_d N_OUT7_Mn8@2467_g N_VSS_Mn8@2467_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2466 N_OUT8_Mn8@2466_d N_OUT7_Mn8@2466_g N_VSS_Mn8@2466_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2467 N_OUT8_Mp8@2467_d N_OUT7_Mp8@2467_g N_VDD_Mp8@2467_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2466 N_OUT8_Mp8@2466_d N_OUT7_Mp8@2466_g N_VDD_Mp8@2466_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2465 N_OUT8_Mn8@2465_d N_OUT7_Mn8@2465_g N_VSS_Mn8@2465_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2464 N_OUT8_Mn8@2464_d N_OUT7_Mn8@2464_g N_VSS_Mn8@2464_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2465 N_OUT8_Mp8@2465_d N_OUT7_Mp8@2465_g N_VDD_Mp8@2465_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2464 N_OUT8_Mp8@2464_d N_OUT7_Mp8@2464_g N_VDD_Mp8@2464_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2463 N_OUT8_Mn8@2463_d N_OUT7_Mn8@2463_g N_VSS_Mn8@2463_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2462 N_OUT8_Mn8@2462_d N_OUT7_Mn8@2462_g N_VSS_Mn8@2462_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2463 N_OUT8_Mp8@2463_d N_OUT7_Mp8@2463_g N_VDD_Mp8@2463_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2462 N_OUT8_Mp8@2462_d N_OUT7_Mp8@2462_g N_VDD_Mp8@2462_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2461 N_OUT8_Mn8@2461_d N_OUT7_Mn8@2461_g N_VSS_Mn8@2461_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2460 N_OUT8_Mn8@2460_d N_OUT7_Mn8@2460_g N_VSS_Mn8@2460_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2461 N_OUT8_Mp8@2461_d N_OUT7_Mp8@2461_g N_VDD_Mp8@2461_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2460 N_OUT8_Mp8@2460_d N_OUT7_Mp8@2460_g N_VDD_Mp8@2460_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2459 N_OUT8_Mn8@2459_d N_OUT7_Mn8@2459_g N_VSS_Mn8@2459_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2458 N_OUT8_Mn8@2458_d N_OUT7_Mn8@2458_g N_VSS_Mn8@2458_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2459 N_OUT8_Mp8@2459_d N_OUT7_Mp8@2459_g N_VDD_Mp8@2459_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2458 N_OUT8_Mp8@2458_d N_OUT7_Mp8@2458_g N_VDD_Mp8@2458_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2457 N_OUT8_Mn8@2457_d N_OUT7_Mn8@2457_g N_VSS_Mn8@2457_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2456 N_OUT8_Mn8@2456_d N_OUT7_Mn8@2456_g N_VSS_Mn8@2456_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2457 N_OUT8_Mp8@2457_d N_OUT7_Mp8@2457_g N_VDD_Mp8@2457_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2456 N_OUT8_Mp8@2456_d N_OUT7_Mp8@2456_g N_VDD_Mp8@2456_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2455 N_OUT8_Mn8@2455_d N_OUT7_Mn8@2455_g N_VSS_Mn8@2455_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2454 N_OUT8_Mn8@2454_d N_OUT7_Mn8@2454_g N_VSS_Mn8@2454_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2455 N_OUT8_Mp8@2455_d N_OUT7_Mp8@2455_g N_VDD_Mp8@2455_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2454 N_OUT8_Mp8@2454_d N_OUT7_Mp8@2454_g N_VDD_Mp8@2454_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2453 N_OUT8_Mn8@2453_d N_OUT7_Mn8@2453_g N_VSS_Mn8@2453_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2452 N_OUT8_Mn8@2452_d N_OUT7_Mn8@2452_g N_VSS_Mn8@2452_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2453 N_OUT8_Mp8@2453_d N_OUT7_Mp8@2453_g N_VDD_Mp8@2453_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2452 N_OUT8_Mp8@2452_d N_OUT7_Mp8@2452_g N_VDD_Mp8@2452_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2451 N_OUT8_Mn8@2451_d N_OUT7_Mn8@2451_g N_VSS_Mn8@2451_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2450 N_OUT8_Mn8@2450_d N_OUT7_Mn8@2450_g N_VSS_Mn8@2450_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2451 N_OUT8_Mp8@2451_d N_OUT7_Mp8@2451_g N_VDD_Mp8@2451_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2450 N_OUT8_Mp8@2450_d N_OUT7_Mp8@2450_g N_VDD_Mp8@2450_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2449 N_OUT8_Mn8@2449_d N_OUT7_Mn8@2449_g N_VSS_Mn8@2449_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2448 N_OUT8_Mn8@2448_d N_OUT7_Mn8@2448_g N_VSS_Mn8@2448_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2449 N_OUT8_Mp8@2449_d N_OUT7_Mp8@2449_g N_VDD_Mp8@2449_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2448 N_OUT8_Mp8@2448_d N_OUT7_Mp8@2448_g N_VDD_Mp8@2448_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2447 N_OUT8_Mn8@2447_d N_OUT7_Mn8@2447_g N_VSS_Mn8@2447_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2446 N_OUT8_Mn8@2446_d N_OUT7_Mn8@2446_g N_VSS_Mn8@2446_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2447 N_OUT8_Mp8@2447_d N_OUT7_Mp8@2447_g N_VDD_Mp8@2447_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2446 N_OUT8_Mp8@2446_d N_OUT7_Mp8@2446_g N_VDD_Mp8@2446_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2445 N_OUT8_Mn8@2445_d N_OUT7_Mn8@2445_g N_VSS_Mn8@2445_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2444 N_OUT8_Mn8@2444_d N_OUT7_Mn8@2444_g N_VSS_Mn8@2444_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2445 N_OUT8_Mp8@2445_d N_OUT7_Mp8@2445_g N_VDD_Mp8@2445_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2444 N_OUT8_Mp8@2444_d N_OUT7_Mp8@2444_g N_VDD_Mp8@2444_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2443 N_OUT8_Mn8@2443_d N_OUT7_Mn8@2443_g N_VSS_Mn8@2443_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2442 N_OUT8_Mn8@2442_d N_OUT7_Mn8@2442_g N_VSS_Mn8@2442_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2443 N_OUT8_Mp8@2443_d N_OUT7_Mp8@2443_g N_VDD_Mp8@2443_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2442 N_OUT8_Mp8@2442_d N_OUT7_Mp8@2442_g N_VDD_Mp8@2442_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2441 N_OUT8_Mn8@2441_d N_OUT7_Mn8@2441_g N_VSS_Mn8@2441_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2440 N_OUT8_Mn8@2440_d N_OUT7_Mn8@2440_g N_VSS_Mn8@2440_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2441 N_OUT8_Mp8@2441_d N_OUT7_Mp8@2441_g N_VDD_Mp8@2441_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2440 N_OUT8_Mp8@2440_d N_OUT7_Mp8@2440_g N_VDD_Mp8@2440_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2439 N_OUT8_Mn8@2439_d N_OUT7_Mn8@2439_g N_VSS_Mn8@2439_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2438 N_OUT8_Mn8@2438_d N_OUT7_Mn8@2438_g N_VSS_Mn8@2438_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2439 N_OUT8_Mp8@2439_d N_OUT7_Mp8@2439_g N_VDD_Mp8@2439_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2438 N_OUT8_Mp8@2438_d N_OUT7_Mp8@2438_g N_VDD_Mp8@2438_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2437 N_OUT8_Mn8@2437_d N_OUT7_Mn8@2437_g N_VSS_Mn8@2437_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2436 N_OUT8_Mn8@2436_d N_OUT7_Mn8@2436_g N_VSS_Mn8@2436_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2437 N_OUT8_Mp8@2437_d N_OUT7_Mp8@2437_g N_VDD_Mp8@2437_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2436 N_OUT8_Mp8@2436_d N_OUT7_Mp8@2436_g N_VDD_Mp8@2436_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2435 N_OUT8_Mn8@2435_d N_OUT7_Mn8@2435_g N_VSS_Mn8@2435_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2434 N_OUT8_Mn8@2434_d N_OUT7_Mn8@2434_g N_VSS_Mn8@2434_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2435 N_OUT8_Mp8@2435_d N_OUT7_Mp8@2435_g N_VDD_Mp8@2435_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2434 N_OUT8_Mp8@2434_d N_OUT7_Mp8@2434_g N_VDD_Mp8@2434_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2433 N_OUT8_Mn8@2433_d N_OUT7_Mn8@2433_g N_VSS_Mn8@2433_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2432 N_OUT8_Mn8@2432_d N_OUT7_Mn8@2432_g N_VSS_Mn8@2432_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2433 N_OUT8_Mp8@2433_d N_OUT7_Mp8@2433_g N_VDD_Mp8@2433_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2432 N_OUT8_Mp8@2432_d N_OUT7_Mp8@2432_g N_VDD_Mp8@2432_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2431 N_OUT8_Mn8@2431_d N_OUT7_Mn8@2431_g N_VSS_Mn8@2431_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2430 N_OUT8_Mn8@2430_d N_OUT7_Mn8@2430_g N_VSS_Mn8@2430_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2431 N_OUT8_Mp8@2431_d N_OUT7_Mp8@2431_g N_VDD_Mp8@2431_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2430 N_OUT8_Mp8@2430_d N_OUT7_Mp8@2430_g N_VDD_Mp8@2430_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2429 N_OUT8_Mn8@2429_d N_OUT7_Mn8@2429_g N_VSS_Mn8@2429_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2428 N_OUT8_Mn8@2428_d N_OUT7_Mn8@2428_g N_VSS_Mn8@2428_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2429 N_OUT8_Mp8@2429_d N_OUT7_Mp8@2429_g N_VDD_Mp8@2429_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2428 N_OUT8_Mp8@2428_d N_OUT7_Mp8@2428_g N_VDD_Mp8@2428_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2427 N_OUT8_Mn8@2427_d N_OUT7_Mn8@2427_g N_VSS_Mn8@2427_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2426 N_OUT8_Mn8@2426_d N_OUT7_Mn8@2426_g N_VSS_Mn8@2426_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2427 N_OUT8_Mp8@2427_d N_OUT7_Mp8@2427_g N_VDD_Mp8@2427_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2426 N_OUT8_Mp8@2426_d N_OUT7_Mp8@2426_g N_VDD_Mp8@2426_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2425 N_OUT8_Mn8@2425_d N_OUT7_Mn8@2425_g N_VSS_Mn8@2425_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2424 N_OUT8_Mn8@2424_d N_OUT7_Mn8@2424_g N_VSS_Mn8@2424_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2425 N_OUT8_Mp8@2425_d N_OUT7_Mp8@2425_g N_VDD_Mp8@2425_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2424 N_OUT8_Mp8@2424_d N_OUT7_Mp8@2424_g N_VDD_Mp8@2424_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2423 N_OUT8_Mn8@2423_d N_OUT7_Mn8@2423_g N_VSS_Mn8@2423_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2422 N_OUT8_Mn8@2422_d N_OUT7_Mn8@2422_g N_VSS_Mn8@2422_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2423 N_OUT8_Mp8@2423_d N_OUT7_Mp8@2423_g N_VDD_Mp8@2423_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2422 N_OUT8_Mp8@2422_d N_OUT7_Mp8@2422_g N_VDD_Mp8@2422_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2421 N_OUT8_Mn8@2421_d N_OUT7_Mn8@2421_g N_VSS_Mn8@2421_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2420 N_OUT8_Mn8@2420_d N_OUT7_Mn8@2420_g N_VSS_Mn8@2420_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2421 N_OUT8_Mp8@2421_d N_OUT7_Mp8@2421_g N_VDD_Mp8@2421_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2420 N_OUT8_Mp8@2420_d N_OUT7_Mp8@2420_g N_VDD_Mp8@2420_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2419 N_OUT8_Mn8@2419_d N_OUT7_Mn8@2419_g N_VSS_Mn8@2419_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2418 N_OUT8_Mn8@2418_d N_OUT7_Mn8@2418_g N_VSS_Mn8@2418_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2419 N_OUT8_Mp8@2419_d N_OUT7_Mp8@2419_g N_VDD_Mp8@2419_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2418 N_OUT8_Mp8@2418_d N_OUT7_Mp8@2418_g N_VDD_Mp8@2418_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2417 N_OUT8_Mn8@2417_d N_OUT7_Mn8@2417_g N_VSS_Mn8@2417_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2416 N_OUT8_Mn8@2416_d N_OUT7_Mn8@2416_g N_VSS_Mn8@2416_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2417 N_OUT8_Mp8@2417_d N_OUT7_Mp8@2417_g N_VDD_Mp8@2417_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2416 N_OUT8_Mp8@2416_d N_OUT7_Mp8@2416_g N_VDD_Mp8@2416_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2415 N_OUT8_Mn8@2415_d N_OUT7_Mn8@2415_g N_VSS_Mn8@2415_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2414 N_OUT8_Mn8@2414_d N_OUT7_Mn8@2414_g N_VSS_Mn8@2414_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2415 N_OUT8_Mp8@2415_d N_OUT7_Mp8@2415_g N_VDD_Mp8@2415_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2414 N_OUT8_Mp8@2414_d N_OUT7_Mp8@2414_g N_VDD_Mp8@2414_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2413 N_OUT8_Mn8@2413_d N_OUT7_Mn8@2413_g N_VSS_Mn8@2413_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2412 N_OUT8_Mn8@2412_d N_OUT7_Mn8@2412_g N_VSS_Mn8@2412_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2413 N_OUT8_Mp8@2413_d N_OUT7_Mp8@2413_g N_VDD_Mp8@2413_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2412 N_OUT8_Mp8@2412_d N_OUT7_Mp8@2412_g N_VDD_Mp8@2412_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2411 N_OUT8_Mn8@2411_d N_OUT7_Mn8@2411_g N_VSS_Mn8@2411_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2410 N_OUT8_Mn8@2410_d N_OUT7_Mn8@2410_g N_VSS_Mn8@2410_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2411 N_OUT8_Mp8@2411_d N_OUT7_Mp8@2411_g N_VDD_Mp8@2411_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2410 N_OUT8_Mp8@2410_d N_OUT7_Mp8@2410_g N_VDD_Mp8@2410_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2409 N_OUT8_Mn8@2409_d N_OUT7_Mn8@2409_g N_VSS_Mn8@2409_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2408 N_OUT8_Mn8@2408_d N_OUT7_Mn8@2408_g N_VSS_Mn8@2408_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2409 N_OUT8_Mp8@2409_d N_OUT7_Mp8@2409_g N_VDD_Mp8@2409_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2408 N_OUT8_Mp8@2408_d N_OUT7_Mp8@2408_g N_VDD_Mp8@2408_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2407 N_OUT8_Mn8@2407_d N_OUT7_Mn8@2407_g N_VSS_Mn8@2407_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2406 N_OUT8_Mn8@2406_d N_OUT7_Mn8@2406_g N_VSS_Mn8@2406_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2407 N_OUT8_Mp8@2407_d N_OUT7_Mp8@2407_g N_VDD_Mp8@2407_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2406 N_OUT8_Mp8@2406_d N_OUT7_Mp8@2406_g N_VDD_Mp8@2406_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2405 N_OUT8_Mn8@2405_d N_OUT7_Mn8@2405_g N_VSS_Mn8@2405_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2404 N_OUT8_Mn8@2404_d N_OUT7_Mn8@2404_g N_VSS_Mn8@2404_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2405 N_OUT8_Mp8@2405_d N_OUT7_Mp8@2405_g N_VDD_Mp8@2405_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2404 N_OUT8_Mp8@2404_d N_OUT7_Mp8@2404_g N_VDD_Mp8@2404_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2403 N_OUT8_Mn8@2403_d N_OUT7_Mn8@2403_g N_VSS_Mn8@2403_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2402 N_OUT8_Mn8@2402_d N_OUT7_Mn8@2402_g N_VSS_Mn8@2402_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2403 N_OUT8_Mp8@2403_d N_OUT7_Mp8@2403_g N_VDD_Mp8@2403_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2402 N_OUT8_Mp8@2402_d N_OUT7_Mp8@2402_g N_VDD_Mp8@2402_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2401 N_OUT8_Mn8@2401_d N_OUT7_Mn8@2401_g N_VSS_Mn8@2401_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2400 N_OUT8_Mn8@2400_d N_OUT7_Mn8@2400_g N_VSS_Mn8@2400_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2401 N_OUT8_Mp8@2401_d N_OUT7_Mp8@2401_g N_VDD_Mp8@2401_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2400 N_OUT8_Mp8@2400_d N_OUT7_Mp8@2400_g N_VDD_Mp8@2400_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2399 N_OUT8_Mn8@2399_d N_OUT7_Mn8@2399_g N_VSS_Mn8@2399_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2398 N_OUT8_Mn8@2398_d N_OUT7_Mn8@2398_g N_VSS_Mn8@2398_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2399 N_OUT8_Mp8@2399_d N_OUT7_Mp8@2399_g N_VDD_Mp8@2399_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2398 N_OUT8_Mp8@2398_d N_OUT7_Mp8@2398_g N_VDD_Mp8@2398_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2397 N_OUT8_Mn8@2397_d N_OUT7_Mn8@2397_g N_VSS_Mn8@2397_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2396 N_OUT8_Mn8@2396_d N_OUT7_Mn8@2396_g N_VSS_Mn8@2396_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2397 N_OUT8_Mp8@2397_d N_OUT7_Mp8@2397_g N_VDD_Mp8@2397_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2396 N_OUT8_Mp8@2396_d N_OUT7_Mp8@2396_g N_VDD_Mp8@2396_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2395 N_OUT8_Mn8@2395_d N_OUT7_Mn8@2395_g N_VSS_Mn8@2395_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2394 N_OUT8_Mn8@2394_d N_OUT7_Mn8@2394_g N_VSS_Mn8@2394_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2395 N_OUT8_Mp8@2395_d N_OUT7_Mp8@2395_g N_VDD_Mp8@2395_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2394 N_OUT8_Mp8@2394_d N_OUT7_Mp8@2394_g N_VDD_Mp8@2394_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2393 N_OUT8_Mn8@2393_d N_OUT7_Mn8@2393_g N_VSS_Mn8@2393_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2392 N_OUT8_Mn8@2392_d N_OUT7_Mn8@2392_g N_VSS_Mn8@2392_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2393 N_OUT8_Mp8@2393_d N_OUT7_Mp8@2393_g N_VDD_Mp8@2393_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2392 N_OUT8_Mp8@2392_d N_OUT7_Mp8@2392_g N_VDD_Mp8@2392_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2391 N_OUT8_Mn8@2391_d N_OUT7_Mn8@2391_g N_VSS_Mn8@2391_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2390 N_OUT8_Mn8@2390_d N_OUT7_Mn8@2390_g N_VSS_Mn8@2390_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2391 N_OUT8_Mp8@2391_d N_OUT7_Mp8@2391_g N_VDD_Mp8@2391_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2390 N_OUT8_Mp8@2390_d N_OUT7_Mp8@2390_g N_VDD_Mp8@2390_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2389 N_OUT8_Mn8@2389_d N_OUT7_Mn8@2389_g N_VSS_Mn8@2389_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2388 N_OUT8_Mn8@2388_d N_OUT7_Mn8@2388_g N_VSS_Mn8@2388_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2389 N_OUT8_Mp8@2389_d N_OUT7_Mp8@2389_g N_VDD_Mp8@2389_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2388 N_OUT8_Mp8@2388_d N_OUT7_Mp8@2388_g N_VDD_Mp8@2388_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2387 N_OUT8_Mn8@2387_d N_OUT7_Mn8@2387_g N_VSS_Mn8@2387_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2386 N_OUT8_Mn8@2386_d N_OUT7_Mn8@2386_g N_VSS_Mn8@2386_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2387 N_OUT8_Mp8@2387_d N_OUT7_Mp8@2387_g N_VDD_Mp8@2387_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2386 N_OUT8_Mp8@2386_d N_OUT7_Mp8@2386_g N_VDD_Mp8@2386_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2385 N_OUT8_Mn8@2385_d N_OUT7_Mn8@2385_g N_VSS_Mn8@2385_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2384 N_OUT8_Mn8@2384_d N_OUT7_Mn8@2384_g N_VSS_Mn8@2384_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2385 N_OUT8_Mp8@2385_d N_OUT7_Mp8@2385_g N_VDD_Mp8@2385_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2384 N_OUT8_Mp8@2384_d N_OUT7_Mp8@2384_g N_VDD_Mp8@2384_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2383 N_OUT8_Mn8@2383_d N_OUT7_Mn8@2383_g N_VSS_Mn8@2383_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2382 N_OUT8_Mn8@2382_d N_OUT7_Mn8@2382_g N_VSS_Mn8@2382_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2383 N_OUT8_Mp8@2383_d N_OUT7_Mp8@2383_g N_VDD_Mp8@2383_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2382 N_OUT8_Mp8@2382_d N_OUT7_Mp8@2382_g N_VDD_Mp8@2382_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2381 N_OUT8_Mn8@2381_d N_OUT7_Mn8@2381_g N_VSS_Mn8@2381_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2380 N_OUT8_Mn8@2380_d N_OUT7_Mn8@2380_g N_VSS_Mn8@2380_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2381 N_OUT8_Mp8@2381_d N_OUT7_Mp8@2381_g N_VDD_Mp8@2381_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2380 N_OUT8_Mp8@2380_d N_OUT7_Mp8@2380_g N_VDD_Mp8@2380_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2379 N_OUT8_Mn8@2379_d N_OUT7_Mn8@2379_g N_VSS_Mn8@2379_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2378 N_OUT8_Mn8@2378_d N_OUT7_Mn8@2378_g N_VSS_Mn8@2378_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2379 N_OUT8_Mp8@2379_d N_OUT7_Mp8@2379_g N_VDD_Mp8@2379_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2378 N_OUT8_Mp8@2378_d N_OUT7_Mp8@2378_g N_VDD_Mp8@2378_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2377 N_OUT8_Mn8@2377_d N_OUT7_Mn8@2377_g N_VSS_Mn8@2377_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2376 N_OUT8_Mn8@2376_d N_OUT7_Mn8@2376_g N_VSS_Mn8@2376_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2377 N_OUT8_Mp8@2377_d N_OUT7_Mp8@2377_g N_VDD_Mp8@2377_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2376 N_OUT8_Mp8@2376_d N_OUT7_Mp8@2376_g N_VDD_Mp8@2376_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2375 N_OUT8_Mn8@2375_d N_OUT7_Mn8@2375_g N_VSS_Mn8@2375_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2374 N_OUT8_Mn8@2374_d N_OUT7_Mn8@2374_g N_VSS_Mn8@2374_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2375 N_OUT8_Mp8@2375_d N_OUT7_Mp8@2375_g N_VDD_Mp8@2375_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2374 N_OUT8_Mp8@2374_d N_OUT7_Mp8@2374_g N_VDD_Mp8@2374_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2373 N_OUT8_Mn8@2373_d N_OUT7_Mn8@2373_g N_VSS_Mn8@2373_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2372 N_OUT8_Mn8@2372_d N_OUT7_Mn8@2372_g N_VSS_Mn8@2372_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2373 N_OUT8_Mp8@2373_d N_OUT7_Mp8@2373_g N_VDD_Mp8@2373_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2372 N_OUT8_Mp8@2372_d N_OUT7_Mp8@2372_g N_VDD_Mp8@2372_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2371 N_OUT8_Mn8@2371_d N_OUT7_Mn8@2371_g N_VSS_Mn8@2371_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2370 N_OUT8_Mn8@2370_d N_OUT7_Mn8@2370_g N_VSS_Mn8@2370_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2371 N_OUT8_Mp8@2371_d N_OUT7_Mp8@2371_g N_VDD_Mp8@2371_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2370 N_OUT8_Mp8@2370_d N_OUT7_Mp8@2370_g N_VDD_Mp8@2370_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2369 N_OUT8_Mn8@2369_d N_OUT7_Mn8@2369_g N_VSS_Mn8@2369_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2368 N_OUT8_Mn8@2368_d N_OUT7_Mn8@2368_g N_VSS_Mn8@2368_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2369 N_OUT8_Mp8@2369_d N_OUT7_Mp8@2369_g N_VDD_Mp8@2369_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2368 N_OUT8_Mp8@2368_d N_OUT7_Mp8@2368_g N_VDD_Mp8@2368_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2367 N_OUT8_Mn8@2367_d N_OUT7_Mn8@2367_g N_VSS_Mn8@2367_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2366 N_OUT8_Mn8@2366_d N_OUT7_Mn8@2366_g N_VSS_Mn8@2366_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2367 N_OUT8_Mp8@2367_d N_OUT7_Mp8@2367_g N_VDD_Mp8@2367_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2366 N_OUT8_Mp8@2366_d N_OUT7_Mp8@2366_g N_VDD_Mp8@2366_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2365 N_OUT8_Mn8@2365_d N_OUT7_Mn8@2365_g N_VSS_Mn8@2365_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2364 N_OUT8_Mn8@2364_d N_OUT7_Mn8@2364_g N_VSS_Mn8@2364_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2365 N_OUT8_Mp8@2365_d N_OUT7_Mp8@2365_g N_VDD_Mp8@2365_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2364 N_OUT8_Mp8@2364_d N_OUT7_Mp8@2364_g N_VDD_Mp8@2364_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2363 N_OUT8_Mn8@2363_d N_OUT7_Mn8@2363_g N_VSS_Mn8@2363_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2362 N_OUT8_Mn8@2362_d N_OUT7_Mn8@2362_g N_VSS_Mn8@2362_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2363 N_OUT8_Mp8@2363_d N_OUT7_Mp8@2363_g N_VDD_Mp8@2363_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2362 N_OUT8_Mp8@2362_d N_OUT7_Mp8@2362_g N_VDD_Mp8@2362_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2361 N_OUT8_Mn8@2361_d N_OUT7_Mn8@2361_g N_VSS_Mn8@2361_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2360 N_OUT8_Mn8@2360_d N_OUT7_Mn8@2360_g N_VSS_Mn8@2360_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2361 N_OUT8_Mp8@2361_d N_OUT7_Mp8@2361_g N_VDD_Mp8@2361_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2360 N_OUT8_Mp8@2360_d N_OUT7_Mp8@2360_g N_VDD_Mp8@2360_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2359 N_OUT8_Mn8@2359_d N_OUT7_Mn8@2359_g N_VSS_Mn8@2359_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2358 N_OUT8_Mn8@2358_d N_OUT7_Mn8@2358_g N_VSS_Mn8@2358_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2359 N_OUT8_Mp8@2359_d N_OUT7_Mp8@2359_g N_VDD_Mp8@2359_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2358 N_OUT8_Mp8@2358_d N_OUT7_Mp8@2358_g N_VDD_Mp8@2358_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2357 N_OUT8_Mn8@2357_d N_OUT7_Mn8@2357_g N_VSS_Mn8@2357_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2356 N_OUT8_Mn8@2356_d N_OUT7_Mn8@2356_g N_VSS_Mn8@2356_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2357 N_OUT8_Mp8@2357_d N_OUT7_Mp8@2357_g N_VDD_Mp8@2357_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2356 N_OUT8_Mp8@2356_d N_OUT7_Mp8@2356_g N_VDD_Mp8@2356_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2355 N_OUT8_Mn8@2355_d N_OUT7_Mn8@2355_g N_VSS_Mn8@2355_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2354 N_OUT8_Mn8@2354_d N_OUT7_Mn8@2354_g N_VSS_Mn8@2354_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2355 N_OUT8_Mp8@2355_d N_OUT7_Mp8@2355_g N_VDD_Mp8@2355_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2354 N_OUT8_Mp8@2354_d N_OUT7_Mp8@2354_g N_VDD_Mp8@2354_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2353 N_OUT8_Mn8@2353_d N_OUT7_Mn8@2353_g N_VSS_Mn8@2353_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2352 N_OUT8_Mn8@2352_d N_OUT7_Mn8@2352_g N_VSS_Mn8@2352_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2353 N_OUT8_Mp8@2353_d N_OUT7_Mp8@2353_g N_VDD_Mp8@2353_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2352 N_OUT8_Mp8@2352_d N_OUT7_Mp8@2352_g N_VDD_Mp8@2352_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2351 N_OUT8_Mn8@2351_d N_OUT7_Mn8@2351_g N_VSS_Mn8@2351_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2350 N_OUT8_Mn8@2350_d N_OUT7_Mn8@2350_g N_VSS_Mn8@2350_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2351 N_OUT8_Mp8@2351_d N_OUT7_Mp8@2351_g N_VDD_Mp8@2351_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2350 N_OUT8_Mp8@2350_d N_OUT7_Mp8@2350_g N_VDD_Mp8@2350_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2349 N_OUT8_Mn8@2349_d N_OUT7_Mn8@2349_g N_VSS_Mn8@2349_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2348 N_OUT8_Mn8@2348_d N_OUT7_Mn8@2348_g N_VSS_Mn8@2348_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2349 N_OUT8_Mp8@2349_d N_OUT7_Mp8@2349_g N_VDD_Mp8@2349_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2348 N_OUT8_Mp8@2348_d N_OUT7_Mp8@2348_g N_VDD_Mp8@2348_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2347 N_OUT8_Mn8@2347_d N_OUT7_Mn8@2347_g N_VSS_Mn8@2347_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2346 N_OUT8_Mn8@2346_d N_OUT7_Mn8@2346_g N_VSS_Mn8@2346_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2347 N_OUT8_Mp8@2347_d N_OUT7_Mp8@2347_g N_VDD_Mp8@2347_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2346 N_OUT8_Mp8@2346_d N_OUT7_Mp8@2346_g N_VDD_Mp8@2346_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2345 N_OUT8_Mn8@2345_d N_OUT7_Mn8@2345_g N_VSS_Mn8@2345_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2344 N_OUT8_Mn8@2344_d N_OUT7_Mn8@2344_g N_VSS_Mn8@2344_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2345 N_OUT8_Mp8@2345_d N_OUT7_Mp8@2345_g N_VDD_Mp8@2345_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2344 N_OUT8_Mp8@2344_d N_OUT7_Mp8@2344_g N_VDD_Mp8@2344_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2343 N_OUT8_Mn8@2343_d N_OUT7_Mn8@2343_g N_VSS_Mn8@2343_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2342 N_OUT8_Mn8@2342_d N_OUT7_Mn8@2342_g N_VSS_Mn8@2342_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2343 N_OUT8_Mp8@2343_d N_OUT7_Mp8@2343_g N_VDD_Mp8@2343_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2342 N_OUT8_Mp8@2342_d N_OUT7_Mp8@2342_g N_VDD_Mp8@2342_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2341 N_OUT8_Mn8@2341_d N_OUT7_Mn8@2341_g N_VSS_Mn8@2341_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2340 N_OUT8_Mn8@2340_d N_OUT7_Mn8@2340_g N_VSS_Mn8@2340_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2341 N_OUT8_Mp8@2341_d N_OUT7_Mp8@2341_g N_VDD_Mp8@2341_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2340 N_OUT8_Mp8@2340_d N_OUT7_Mp8@2340_g N_VDD_Mp8@2340_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2339 N_OUT8_Mn8@2339_d N_OUT7_Mn8@2339_g N_VSS_Mn8@2339_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2338 N_OUT8_Mn8@2338_d N_OUT7_Mn8@2338_g N_VSS_Mn8@2338_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2339 N_OUT8_Mp8@2339_d N_OUT7_Mp8@2339_g N_VDD_Mp8@2339_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2338 N_OUT8_Mp8@2338_d N_OUT7_Mp8@2338_g N_VDD_Mp8@2338_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2337 N_OUT8_Mn8@2337_d N_OUT7_Mn8@2337_g N_VSS_Mn8@2337_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2336 N_OUT8_Mn8@2336_d N_OUT7_Mn8@2336_g N_VSS_Mn8@2336_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2337 N_OUT8_Mp8@2337_d N_OUT7_Mp8@2337_g N_VDD_Mp8@2337_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2336 N_OUT8_Mp8@2336_d N_OUT7_Mp8@2336_g N_VDD_Mp8@2336_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2335 N_OUT8_Mn8@2335_d N_OUT7_Mn8@2335_g N_VSS_Mn8@2335_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2334 N_OUT8_Mn8@2334_d N_OUT7_Mn8@2334_g N_VSS_Mn8@2334_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2335 N_OUT8_Mp8@2335_d N_OUT7_Mp8@2335_g N_VDD_Mp8@2335_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2334 N_OUT8_Mp8@2334_d N_OUT7_Mp8@2334_g N_VDD_Mp8@2334_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2333 N_OUT8_Mn8@2333_d N_OUT7_Mn8@2333_g N_VSS_Mn8@2333_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2332 N_OUT8_Mn8@2332_d N_OUT7_Mn8@2332_g N_VSS_Mn8@2332_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2333 N_OUT8_Mp8@2333_d N_OUT7_Mp8@2333_g N_VDD_Mp8@2333_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2332 N_OUT8_Mp8@2332_d N_OUT7_Mp8@2332_g N_VDD_Mp8@2332_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2331 N_OUT8_Mn8@2331_d N_OUT7_Mn8@2331_g N_VSS_Mn8@2331_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2330 N_OUT8_Mn8@2330_d N_OUT7_Mn8@2330_g N_VSS_Mn8@2330_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2331 N_OUT8_Mp8@2331_d N_OUT7_Mp8@2331_g N_VDD_Mp8@2331_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2330 N_OUT8_Mp8@2330_d N_OUT7_Mp8@2330_g N_VDD_Mp8@2330_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2329 N_OUT8_Mn8@2329_d N_OUT7_Mn8@2329_g N_VSS_Mn8@2329_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2328 N_OUT8_Mn8@2328_d N_OUT7_Mn8@2328_g N_VSS_Mn8@2328_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2329 N_OUT8_Mp8@2329_d N_OUT7_Mp8@2329_g N_VDD_Mp8@2329_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2328 N_OUT8_Mp8@2328_d N_OUT7_Mp8@2328_g N_VDD_Mp8@2328_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2327 N_OUT8_Mn8@2327_d N_OUT7_Mn8@2327_g N_VSS_Mn8@2327_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2326 N_OUT8_Mn8@2326_d N_OUT7_Mn8@2326_g N_VSS_Mn8@2326_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2327 N_OUT8_Mp8@2327_d N_OUT7_Mp8@2327_g N_VDD_Mp8@2327_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2326 N_OUT8_Mp8@2326_d N_OUT7_Mp8@2326_g N_VDD_Mp8@2326_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2325 N_OUT8_Mn8@2325_d N_OUT7_Mn8@2325_g N_VSS_Mn8@2325_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2324 N_OUT8_Mn8@2324_d N_OUT7_Mn8@2324_g N_VSS_Mn8@2324_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2325 N_OUT8_Mp8@2325_d N_OUT7_Mp8@2325_g N_VDD_Mp8@2325_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2324 N_OUT8_Mp8@2324_d N_OUT7_Mp8@2324_g N_VDD_Mp8@2324_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2323 N_OUT8_Mn8@2323_d N_OUT7_Mn8@2323_g N_VSS_Mn8@2323_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2322 N_OUT8_Mn8@2322_d N_OUT7_Mn8@2322_g N_VSS_Mn8@2322_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2323 N_OUT8_Mp8@2323_d N_OUT7_Mp8@2323_g N_VDD_Mp8@2323_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2322 N_OUT8_Mp8@2322_d N_OUT7_Mp8@2322_g N_VDD_Mp8@2322_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2321 N_OUT8_Mn8@2321_d N_OUT7_Mn8@2321_g N_VSS_Mn8@2321_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2320 N_OUT8_Mn8@2320_d N_OUT7_Mn8@2320_g N_VSS_Mn8@2320_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2321 N_OUT8_Mp8@2321_d N_OUT7_Mp8@2321_g N_VDD_Mp8@2321_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2320 N_OUT8_Mp8@2320_d N_OUT7_Mp8@2320_g N_VDD_Mp8@2320_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2319 N_OUT8_Mn8@2319_d N_OUT7_Mn8@2319_g N_VSS_Mn8@2319_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2318 N_OUT8_Mn8@2318_d N_OUT7_Mn8@2318_g N_VSS_Mn8@2318_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2319 N_OUT8_Mp8@2319_d N_OUT7_Mp8@2319_g N_VDD_Mp8@2319_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2318 N_OUT8_Mp8@2318_d N_OUT7_Mp8@2318_g N_VDD_Mp8@2318_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2317 N_OUT8_Mn8@2317_d N_OUT7_Mn8@2317_g N_VSS_Mn8@2317_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2316 N_OUT8_Mn8@2316_d N_OUT7_Mn8@2316_g N_VSS_Mn8@2316_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2317 N_OUT8_Mp8@2317_d N_OUT7_Mp8@2317_g N_VDD_Mp8@2317_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2316 N_OUT8_Mp8@2316_d N_OUT7_Mp8@2316_g N_VDD_Mp8@2316_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2315 N_OUT8_Mn8@2315_d N_OUT7_Mn8@2315_g N_VSS_Mn8@2315_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2314 N_OUT8_Mn8@2314_d N_OUT7_Mn8@2314_g N_VSS_Mn8@2314_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2315 N_OUT8_Mp8@2315_d N_OUT7_Mp8@2315_g N_VDD_Mp8@2315_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2314 N_OUT8_Mp8@2314_d N_OUT7_Mp8@2314_g N_VDD_Mp8@2314_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2313 N_OUT8_Mn8@2313_d N_OUT7_Mn8@2313_g N_VSS_Mn8@2313_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2312 N_OUT8_Mn8@2312_d N_OUT7_Mn8@2312_g N_VSS_Mn8@2312_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2313 N_OUT8_Mp8@2313_d N_OUT7_Mp8@2313_g N_VDD_Mp8@2313_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2312 N_OUT8_Mp8@2312_d N_OUT7_Mp8@2312_g N_VDD_Mp8@2312_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2311 N_OUT8_Mn8@2311_d N_OUT7_Mn8@2311_g N_VSS_Mn8@2311_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2310 N_OUT8_Mn8@2310_d N_OUT7_Mn8@2310_g N_VSS_Mn8@2310_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2311 N_OUT8_Mp8@2311_d N_OUT7_Mp8@2311_g N_VDD_Mp8@2311_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2310 N_OUT8_Mp8@2310_d N_OUT7_Mp8@2310_g N_VDD_Mp8@2310_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2309 N_OUT8_Mn8@2309_d N_OUT7_Mn8@2309_g N_VSS_Mn8@2309_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2308 N_OUT8_Mn8@2308_d N_OUT7_Mn8@2308_g N_VSS_Mn8@2308_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2309 N_OUT8_Mp8@2309_d N_OUT7_Mp8@2309_g N_VDD_Mp8@2309_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2308 N_OUT8_Mp8@2308_d N_OUT7_Mp8@2308_g N_VDD_Mp8@2308_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2307 N_OUT8_Mn8@2307_d N_OUT7_Mn8@2307_g N_VSS_Mn8@2307_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2306 N_OUT8_Mn8@2306_d N_OUT7_Mn8@2306_g N_VSS_Mn8@2306_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2307 N_OUT8_Mp8@2307_d N_OUT7_Mp8@2307_g N_VDD_Mp8@2307_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2306 N_OUT8_Mp8@2306_d N_OUT7_Mp8@2306_g N_VDD_Mp8@2306_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2305 N_OUT8_Mn8@2305_d N_OUT7_Mn8@2305_g N_VSS_Mn8@2305_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2304 N_OUT8_Mn8@2304_d N_OUT7_Mn8@2304_g N_VSS_Mn8@2304_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2305 N_OUT8_Mp8@2305_d N_OUT7_Mp8@2305_g N_VDD_Mp8@2305_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2304 N_OUT8_Mp8@2304_d N_OUT7_Mp8@2304_g N_VDD_Mp8@2304_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2303 N_OUT8_Mn8@2303_d N_OUT7_Mn8@2303_g N_VSS_Mn8@2303_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2302 N_OUT8_Mn8@2302_d N_OUT7_Mn8@2302_g N_VSS_Mn8@2302_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2303 N_OUT8_Mp8@2303_d N_OUT7_Mp8@2303_g N_VDD_Mp8@2303_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2302 N_OUT8_Mp8@2302_d N_OUT7_Mp8@2302_g N_VDD_Mp8@2302_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2301 N_OUT8_Mn8@2301_d N_OUT7_Mn8@2301_g N_VSS_Mn8@2301_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2300 N_OUT8_Mn8@2300_d N_OUT7_Mn8@2300_g N_VSS_Mn8@2300_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2301 N_OUT8_Mp8@2301_d N_OUT7_Mp8@2301_g N_VDD_Mp8@2301_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2300 N_OUT8_Mp8@2300_d N_OUT7_Mp8@2300_g N_VDD_Mp8@2300_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2299 N_OUT8_Mn8@2299_d N_OUT7_Mn8@2299_g N_VSS_Mn8@2299_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2298 N_OUT8_Mn8@2298_d N_OUT7_Mn8@2298_g N_VSS_Mn8@2298_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2299 N_OUT8_Mp8@2299_d N_OUT7_Mp8@2299_g N_VDD_Mp8@2299_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2298 N_OUT8_Mp8@2298_d N_OUT7_Mp8@2298_g N_VDD_Mp8@2298_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2297 N_OUT8_Mn8@2297_d N_OUT7_Mn8@2297_g N_VSS_Mn8@2297_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2296 N_OUT8_Mn8@2296_d N_OUT7_Mn8@2296_g N_VSS_Mn8@2296_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2297 N_OUT8_Mp8@2297_d N_OUT7_Mp8@2297_g N_VDD_Mp8@2297_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2296 N_OUT8_Mp8@2296_d N_OUT7_Mp8@2296_g N_VDD_Mp8@2296_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2295 N_OUT8_Mn8@2295_d N_OUT7_Mn8@2295_g N_VSS_Mn8@2295_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2294 N_OUT8_Mn8@2294_d N_OUT7_Mn8@2294_g N_VSS_Mn8@2294_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2295 N_OUT8_Mp8@2295_d N_OUT7_Mp8@2295_g N_VDD_Mp8@2295_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2294 N_OUT8_Mp8@2294_d N_OUT7_Mp8@2294_g N_VDD_Mp8@2294_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2293 N_OUT8_Mn8@2293_d N_OUT7_Mn8@2293_g N_VSS_Mn8@2293_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2292 N_OUT8_Mn8@2292_d N_OUT7_Mn8@2292_g N_VSS_Mn8@2292_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2293 N_OUT8_Mp8@2293_d N_OUT7_Mp8@2293_g N_VDD_Mp8@2293_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2292 N_OUT8_Mp8@2292_d N_OUT7_Mp8@2292_g N_VDD_Mp8@2292_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2291 N_OUT8_Mn8@2291_d N_OUT7_Mn8@2291_g N_VSS_Mn8@2291_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2290 N_OUT8_Mn8@2290_d N_OUT7_Mn8@2290_g N_VSS_Mn8@2290_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2291 N_OUT8_Mp8@2291_d N_OUT7_Mp8@2291_g N_VDD_Mp8@2291_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2290 N_OUT8_Mp8@2290_d N_OUT7_Mp8@2290_g N_VDD_Mp8@2290_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2289 N_OUT8_Mn8@2289_d N_OUT7_Mn8@2289_g N_VSS_Mn8@2289_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2288 N_OUT8_Mn8@2288_d N_OUT7_Mn8@2288_g N_VSS_Mn8@2288_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2289 N_OUT8_Mp8@2289_d N_OUT7_Mp8@2289_g N_VDD_Mp8@2289_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2288 N_OUT8_Mp8@2288_d N_OUT7_Mp8@2288_g N_VDD_Mp8@2288_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2287 N_OUT8_Mn8@2287_d N_OUT7_Mn8@2287_g N_VSS_Mn8@2287_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2286 N_OUT8_Mn8@2286_d N_OUT7_Mn8@2286_g N_VSS_Mn8@2286_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2287 N_OUT8_Mp8@2287_d N_OUT7_Mp8@2287_g N_VDD_Mp8@2287_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2286 N_OUT8_Mp8@2286_d N_OUT7_Mp8@2286_g N_VDD_Mp8@2286_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2285 N_OUT8_Mn8@2285_d N_OUT7_Mn8@2285_g N_VSS_Mn8@2285_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2284 N_OUT8_Mn8@2284_d N_OUT7_Mn8@2284_g N_VSS_Mn8@2284_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2285 N_OUT8_Mp8@2285_d N_OUT7_Mp8@2285_g N_VDD_Mp8@2285_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2284 N_OUT8_Mp8@2284_d N_OUT7_Mp8@2284_g N_VDD_Mp8@2284_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2283 N_OUT8_Mn8@2283_d N_OUT7_Mn8@2283_g N_VSS_Mn8@2283_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2282 N_OUT8_Mn8@2282_d N_OUT7_Mn8@2282_g N_VSS_Mn8@2282_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2283 N_OUT8_Mp8@2283_d N_OUT7_Mp8@2283_g N_VDD_Mp8@2283_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2282 N_OUT8_Mp8@2282_d N_OUT7_Mp8@2282_g N_VDD_Mp8@2282_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2281 N_OUT8_Mn8@2281_d N_OUT7_Mn8@2281_g N_VSS_Mn8@2281_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2280 N_OUT8_Mn8@2280_d N_OUT7_Mn8@2280_g N_VSS_Mn8@2280_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2281 N_OUT8_Mp8@2281_d N_OUT7_Mp8@2281_g N_VDD_Mp8@2281_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2280 N_OUT8_Mp8@2280_d N_OUT7_Mp8@2280_g N_VDD_Mp8@2280_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2279 N_OUT8_Mn8@2279_d N_OUT7_Mn8@2279_g N_VSS_Mn8@2279_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2278 N_OUT8_Mn8@2278_d N_OUT7_Mn8@2278_g N_VSS_Mn8@2278_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2279 N_OUT8_Mp8@2279_d N_OUT7_Mp8@2279_g N_VDD_Mp8@2279_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2278 N_OUT8_Mp8@2278_d N_OUT7_Mp8@2278_g N_VDD_Mp8@2278_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2277 N_OUT8_Mn8@2277_d N_OUT7_Mn8@2277_g N_VSS_Mn8@2277_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2276 N_OUT8_Mn8@2276_d N_OUT7_Mn8@2276_g N_VSS_Mn8@2276_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2277 N_OUT8_Mp8@2277_d N_OUT7_Mp8@2277_g N_VDD_Mp8@2277_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2276 N_OUT8_Mp8@2276_d N_OUT7_Mp8@2276_g N_VDD_Mp8@2276_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2275 N_OUT8_Mn8@2275_d N_OUT7_Mn8@2275_g N_VSS_Mn8@2275_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2274 N_OUT8_Mn8@2274_d N_OUT7_Mn8@2274_g N_VSS_Mn8@2274_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2275 N_OUT8_Mp8@2275_d N_OUT7_Mp8@2275_g N_VDD_Mp8@2275_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2274 N_OUT8_Mp8@2274_d N_OUT7_Mp8@2274_g N_VDD_Mp8@2274_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2273 N_OUT8_Mn8@2273_d N_OUT7_Mn8@2273_g N_VSS_Mn8@2273_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2272 N_OUT8_Mn8@2272_d N_OUT7_Mn8@2272_g N_VSS_Mn8@2272_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2273 N_OUT8_Mp8@2273_d N_OUT7_Mp8@2273_g N_VDD_Mp8@2273_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2272 N_OUT8_Mp8@2272_d N_OUT7_Mp8@2272_g N_VDD_Mp8@2272_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2271 N_OUT8_Mn8@2271_d N_OUT7_Mn8@2271_g N_VSS_Mn8@2271_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2270 N_OUT8_Mn8@2270_d N_OUT7_Mn8@2270_g N_VSS_Mn8@2270_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2271 N_OUT8_Mp8@2271_d N_OUT7_Mp8@2271_g N_VDD_Mp8@2271_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2270 N_OUT8_Mp8@2270_d N_OUT7_Mp8@2270_g N_VDD_Mp8@2270_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2269 N_OUT8_Mn8@2269_d N_OUT7_Mn8@2269_g N_VSS_Mn8@2269_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2268 N_OUT8_Mn8@2268_d N_OUT7_Mn8@2268_g N_VSS_Mn8@2268_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2269 N_OUT8_Mp8@2269_d N_OUT7_Mp8@2269_g N_VDD_Mp8@2269_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2268 N_OUT8_Mp8@2268_d N_OUT7_Mp8@2268_g N_VDD_Mp8@2268_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2267 N_OUT8_Mn8@2267_d N_OUT7_Mn8@2267_g N_VSS_Mn8@2267_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2266 N_OUT8_Mn8@2266_d N_OUT7_Mn8@2266_g N_VSS_Mn8@2266_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2267 N_OUT8_Mp8@2267_d N_OUT7_Mp8@2267_g N_VDD_Mp8@2267_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2266 N_OUT8_Mp8@2266_d N_OUT7_Mp8@2266_g N_VDD_Mp8@2266_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2265 N_OUT8_Mn8@2265_d N_OUT7_Mn8@2265_g N_VSS_Mn8@2265_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2264 N_OUT8_Mn8@2264_d N_OUT7_Mn8@2264_g N_VSS_Mn8@2264_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2265 N_OUT8_Mp8@2265_d N_OUT7_Mp8@2265_g N_VDD_Mp8@2265_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2264 N_OUT8_Mp8@2264_d N_OUT7_Mp8@2264_g N_VDD_Mp8@2264_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2263 N_OUT8_Mn8@2263_d N_OUT7_Mn8@2263_g N_VSS_Mn8@2263_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2262 N_OUT8_Mn8@2262_d N_OUT7_Mn8@2262_g N_VSS_Mn8@2262_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2263 N_OUT8_Mp8@2263_d N_OUT7_Mp8@2263_g N_VDD_Mp8@2263_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2262 N_OUT8_Mp8@2262_d N_OUT7_Mp8@2262_g N_VDD_Mp8@2262_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2261 N_OUT8_Mn8@2261_d N_OUT7_Mn8@2261_g N_VSS_Mn8@2261_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2260 N_OUT8_Mn8@2260_d N_OUT7_Mn8@2260_g N_VSS_Mn8@2260_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2261 N_OUT8_Mp8@2261_d N_OUT7_Mp8@2261_g N_VDD_Mp8@2261_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2260 N_OUT8_Mp8@2260_d N_OUT7_Mp8@2260_g N_VDD_Mp8@2260_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2259 N_OUT8_Mn8@2259_d N_OUT7_Mn8@2259_g N_VSS_Mn8@2259_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2258 N_OUT8_Mn8@2258_d N_OUT7_Mn8@2258_g N_VSS_Mn8@2258_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2259 N_OUT8_Mp8@2259_d N_OUT7_Mp8@2259_g N_VDD_Mp8@2259_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2258 N_OUT8_Mp8@2258_d N_OUT7_Mp8@2258_g N_VDD_Mp8@2258_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2257 N_OUT8_Mn8@2257_d N_OUT7_Mn8@2257_g N_VSS_Mn8@2257_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2256 N_OUT8_Mn8@2256_d N_OUT7_Mn8@2256_g N_VSS_Mn8@2256_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2257 N_OUT8_Mp8@2257_d N_OUT7_Mp8@2257_g N_VDD_Mp8@2257_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2256 N_OUT8_Mp8@2256_d N_OUT7_Mp8@2256_g N_VDD_Mp8@2256_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2255 N_OUT8_Mn8@2255_d N_OUT7_Mn8@2255_g N_VSS_Mn8@2255_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2254 N_OUT8_Mn8@2254_d N_OUT7_Mn8@2254_g N_VSS_Mn8@2254_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2255 N_OUT8_Mp8@2255_d N_OUT7_Mp8@2255_g N_VDD_Mp8@2255_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2254 N_OUT8_Mp8@2254_d N_OUT7_Mp8@2254_g N_VDD_Mp8@2254_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2253 N_OUT8_Mn8@2253_d N_OUT7_Mn8@2253_g N_VSS_Mn8@2253_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2252 N_OUT8_Mn8@2252_d N_OUT7_Mn8@2252_g N_VSS_Mn8@2252_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2253 N_OUT8_Mp8@2253_d N_OUT7_Mp8@2253_g N_VDD_Mp8@2253_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2252 N_OUT8_Mp8@2252_d N_OUT7_Mp8@2252_g N_VDD_Mp8@2252_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2251 N_OUT8_Mn8@2251_d N_OUT7_Mn8@2251_g N_VSS_Mn8@2251_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2250 N_OUT8_Mn8@2250_d N_OUT7_Mn8@2250_g N_VSS_Mn8@2250_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2251 N_OUT8_Mp8@2251_d N_OUT7_Mp8@2251_g N_VDD_Mp8@2251_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2250 N_OUT8_Mp8@2250_d N_OUT7_Mp8@2250_g N_VDD_Mp8@2250_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2249 N_OUT8_Mn8@2249_d N_OUT7_Mn8@2249_g N_VSS_Mn8@2249_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2248 N_OUT8_Mn8@2248_d N_OUT7_Mn8@2248_g N_VSS_Mn8@2248_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2249 N_OUT8_Mp8@2249_d N_OUT7_Mp8@2249_g N_VDD_Mp8@2249_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2248 N_OUT8_Mp8@2248_d N_OUT7_Mp8@2248_g N_VDD_Mp8@2248_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2247 N_OUT8_Mn8@2247_d N_OUT7_Mn8@2247_g N_VSS_Mn8@2247_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2246 N_OUT8_Mn8@2246_d N_OUT7_Mn8@2246_g N_VSS_Mn8@2246_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2247 N_OUT8_Mp8@2247_d N_OUT7_Mp8@2247_g N_VDD_Mp8@2247_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2246 N_OUT8_Mp8@2246_d N_OUT7_Mp8@2246_g N_VDD_Mp8@2246_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2245 N_OUT8_Mn8@2245_d N_OUT7_Mn8@2245_g N_VSS_Mn8@2245_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2244 N_OUT8_Mn8@2244_d N_OUT7_Mn8@2244_g N_VSS_Mn8@2244_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2245 N_OUT8_Mp8@2245_d N_OUT7_Mp8@2245_g N_VDD_Mp8@2245_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2244 N_OUT8_Mp8@2244_d N_OUT7_Mp8@2244_g N_VDD_Mp8@2244_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2243 N_OUT8_Mn8@2243_d N_OUT7_Mn8@2243_g N_VSS_Mn8@2243_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2242 N_OUT8_Mn8@2242_d N_OUT7_Mn8@2242_g N_VSS_Mn8@2242_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2243 N_OUT8_Mp8@2243_d N_OUT7_Mp8@2243_g N_VDD_Mp8@2243_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2242 N_OUT8_Mp8@2242_d N_OUT7_Mp8@2242_g N_VDD_Mp8@2242_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2241 N_OUT8_Mn8@2241_d N_OUT7_Mn8@2241_g N_VSS_Mn8@2241_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2240 N_OUT8_Mn8@2240_d N_OUT7_Mn8@2240_g N_VSS_Mn8@2240_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2241 N_OUT8_Mp8@2241_d N_OUT7_Mp8@2241_g N_VDD_Mp8@2241_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2240 N_OUT8_Mp8@2240_d N_OUT7_Mp8@2240_g N_VDD_Mp8@2240_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2239 N_OUT8_Mn8@2239_d N_OUT7_Mn8@2239_g N_VSS_Mn8@2239_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2238 N_OUT8_Mn8@2238_d N_OUT7_Mn8@2238_g N_VSS_Mn8@2238_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2239 N_OUT8_Mp8@2239_d N_OUT7_Mp8@2239_g N_VDD_Mp8@2239_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2238 N_OUT8_Mp8@2238_d N_OUT7_Mp8@2238_g N_VDD_Mp8@2238_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2237 N_OUT8_Mn8@2237_d N_OUT7_Mn8@2237_g N_VSS_Mn8@2237_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2236 N_OUT8_Mn8@2236_d N_OUT7_Mn8@2236_g N_VSS_Mn8@2236_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2237 N_OUT8_Mp8@2237_d N_OUT7_Mp8@2237_g N_VDD_Mp8@2237_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2236 N_OUT8_Mp8@2236_d N_OUT7_Mp8@2236_g N_VDD_Mp8@2236_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2235 N_OUT8_Mn8@2235_d N_OUT7_Mn8@2235_g N_VSS_Mn8@2235_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2234 N_OUT8_Mn8@2234_d N_OUT7_Mn8@2234_g N_VSS_Mn8@2234_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2235 N_OUT8_Mp8@2235_d N_OUT7_Mp8@2235_g N_VDD_Mp8@2235_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2234 N_OUT8_Mp8@2234_d N_OUT7_Mp8@2234_g N_VDD_Mp8@2234_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2233 N_OUT8_Mn8@2233_d N_OUT7_Mn8@2233_g N_VSS_Mn8@2233_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2232 N_OUT8_Mn8@2232_d N_OUT7_Mn8@2232_g N_VSS_Mn8@2232_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2233 N_OUT8_Mp8@2233_d N_OUT7_Mp8@2233_g N_VDD_Mp8@2233_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2232 N_OUT8_Mp8@2232_d N_OUT7_Mp8@2232_g N_VDD_Mp8@2232_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2231 N_OUT8_Mn8@2231_d N_OUT7_Mn8@2231_g N_VSS_Mn8@2231_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2230 N_OUT8_Mn8@2230_d N_OUT7_Mn8@2230_g N_VSS_Mn8@2230_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2231 N_OUT8_Mp8@2231_d N_OUT7_Mp8@2231_g N_VDD_Mp8@2231_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2230 N_OUT8_Mp8@2230_d N_OUT7_Mp8@2230_g N_VDD_Mp8@2230_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2229 N_OUT8_Mn8@2229_d N_OUT7_Mn8@2229_g N_VSS_Mn8@2229_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2228 N_OUT8_Mn8@2228_d N_OUT7_Mn8@2228_g N_VSS_Mn8@2228_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2229 N_OUT8_Mp8@2229_d N_OUT7_Mp8@2229_g N_VDD_Mp8@2229_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2228 N_OUT8_Mp8@2228_d N_OUT7_Mp8@2228_g N_VDD_Mp8@2228_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2227 N_OUT8_Mn8@2227_d N_OUT7_Mn8@2227_g N_VSS_Mn8@2227_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2226 N_OUT8_Mn8@2226_d N_OUT7_Mn8@2226_g N_VSS_Mn8@2226_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2227 N_OUT8_Mp8@2227_d N_OUT7_Mp8@2227_g N_VDD_Mp8@2227_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2226 N_OUT8_Mp8@2226_d N_OUT7_Mp8@2226_g N_VDD_Mp8@2226_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2225 N_OUT8_Mn8@2225_d N_OUT7_Mn8@2225_g N_VSS_Mn8@2225_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2224 N_OUT8_Mn8@2224_d N_OUT7_Mn8@2224_g N_VSS_Mn8@2224_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2225 N_OUT8_Mp8@2225_d N_OUT7_Mp8@2225_g N_VDD_Mp8@2225_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2224 N_OUT8_Mp8@2224_d N_OUT7_Mp8@2224_g N_VDD_Mp8@2224_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2223 N_OUT8_Mn8@2223_d N_OUT7_Mn8@2223_g N_VSS_Mn8@2223_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2222 N_OUT8_Mn8@2222_d N_OUT7_Mn8@2222_g N_VSS_Mn8@2222_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2223 N_OUT8_Mp8@2223_d N_OUT7_Mp8@2223_g N_VDD_Mp8@2223_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2222 N_OUT8_Mp8@2222_d N_OUT7_Mp8@2222_g N_VDD_Mp8@2222_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2221 N_OUT8_Mn8@2221_d N_OUT7_Mn8@2221_g N_VSS_Mn8@2221_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2220 N_OUT8_Mn8@2220_d N_OUT7_Mn8@2220_g N_VSS_Mn8@2220_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2221 N_OUT8_Mp8@2221_d N_OUT7_Mp8@2221_g N_VDD_Mp8@2221_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2220 N_OUT8_Mp8@2220_d N_OUT7_Mp8@2220_g N_VDD_Mp8@2220_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2219 N_OUT8_Mn8@2219_d N_OUT7_Mn8@2219_g N_VSS_Mn8@2219_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2218 N_OUT8_Mn8@2218_d N_OUT7_Mn8@2218_g N_VSS_Mn8@2218_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2219 N_OUT8_Mp8@2219_d N_OUT7_Mp8@2219_g N_VDD_Mp8@2219_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2218 N_OUT8_Mp8@2218_d N_OUT7_Mp8@2218_g N_VDD_Mp8@2218_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2217 N_OUT8_Mn8@2217_d N_OUT7_Mn8@2217_g N_VSS_Mn8@2217_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2216 N_OUT8_Mn8@2216_d N_OUT7_Mn8@2216_g N_VSS_Mn8@2216_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2217 N_OUT8_Mp8@2217_d N_OUT7_Mp8@2217_g N_VDD_Mp8@2217_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2216 N_OUT8_Mp8@2216_d N_OUT7_Mp8@2216_g N_VDD_Mp8@2216_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2215 N_OUT8_Mn8@2215_d N_OUT7_Mn8@2215_g N_VSS_Mn8@2215_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2214 N_OUT8_Mn8@2214_d N_OUT7_Mn8@2214_g N_VSS_Mn8@2214_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2215 N_OUT8_Mp8@2215_d N_OUT7_Mp8@2215_g N_VDD_Mp8@2215_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2214 N_OUT8_Mp8@2214_d N_OUT7_Mp8@2214_g N_VDD_Mp8@2214_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2213 N_OUT8_Mn8@2213_d N_OUT7_Mn8@2213_g N_VSS_Mn8@2213_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2212 N_OUT8_Mn8@2212_d N_OUT7_Mn8@2212_g N_VSS_Mn8@2212_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2213 N_OUT8_Mp8@2213_d N_OUT7_Mp8@2213_g N_VDD_Mp8@2213_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2212 N_OUT8_Mp8@2212_d N_OUT7_Mp8@2212_g N_VDD_Mp8@2212_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2211 N_OUT8_Mn8@2211_d N_OUT7_Mn8@2211_g N_VSS_Mn8@2211_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2210 N_OUT8_Mn8@2210_d N_OUT7_Mn8@2210_g N_VSS_Mn8@2210_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2211 N_OUT8_Mp8@2211_d N_OUT7_Mp8@2211_g N_VDD_Mp8@2211_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2210 N_OUT8_Mp8@2210_d N_OUT7_Mp8@2210_g N_VDD_Mp8@2210_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2209 N_OUT8_Mn8@2209_d N_OUT7_Mn8@2209_g N_VSS_Mn8@2209_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2208 N_OUT8_Mn8@2208_d N_OUT7_Mn8@2208_g N_VSS_Mn8@2208_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2209 N_OUT8_Mp8@2209_d N_OUT7_Mp8@2209_g N_VDD_Mp8@2209_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2208 N_OUT8_Mp8@2208_d N_OUT7_Mp8@2208_g N_VDD_Mp8@2208_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2207 N_OUT8_Mn8@2207_d N_OUT7_Mn8@2207_g N_VSS_Mn8@2207_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2206 N_OUT8_Mn8@2206_d N_OUT7_Mn8@2206_g N_VSS_Mn8@2206_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2207 N_OUT8_Mp8@2207_d N_OUT7_Mp8@2207_g N_VDD_Mp8@2207_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2206 N_OUT8_Mp8@2206_d N_OUT7_Mp8@2206_g N_VDD_Mp8@2206_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2205 N_OUT8_Mn8@2205_d N_OUT7_Mn8@2205_g N_VSS_Mn8@2205_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2204 N_OUT8_Mn8@2204_d N_OUT7_Mn8@2204_g N_VSS_Mn8@2204_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2205 N_OUT8_Mp8@2205_d N_OUT7_Mp8@2205_g N_VDD_Mp8@2205_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2204 N_OUT8_Mp8@2204_d N_OUT7_Mp8@2204_g N_VDD_Mp8@2204_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2203 N_OUT8_Mn8@2203_d N_OUT7_Mn8@2203_g N_VSS_Mn8@2203_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2202 N_OUT8_Mn8@2202_d N_OUT7_Mn8@2202_g N_VSS_Mn8@2202_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2203 N_OUT8_Mp8@2203_d N_OUT7_Mp8@2203_g N_VDD_Mp8@2203_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2202 N_OUT8_Mp8@2202_d N_OUT7_Mp8@2202_g N_VDD_Mp8@2202_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2201 N_OUT8_Mn8@2201_d N_OUT7_Mn8@2201_g N_VSS_Mn8@2201_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2200 N_OUT8_Mn8@2200_d N_OUT7_Mn8@2200_g N_VSS_Mn8@2200_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2201 N_OUT8_Mp8@2201_d N_OUT7_Mp8@2201_g N_VDD_Mp8@2201_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2200 N_OUT8_Mp8@2200_d N_OUT7_Mp8@2200_g N_VDD_Mp8@2200_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2199 N_OUT8_Mn8@2199_d N_OUT7_Mn8@2199_g N_VSS_Mn8@2199_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2198 N_OUT8_Mn8@2198_d N_OUT7_Mn8@2198_g N_VSS_Mn8@2198_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2199 N_OUT8_Mp8@2199_d N_OUT7_Mp8@2199_g N_VDD_Mp8@2199_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2198 N_OUT8_Mp8@2198_d N_OUT7_Mp8@2198_g N_VDD_Mp8@2198_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2197 N_OUT8_Mn8@2197_d N_OUT7_Mn8@2197_g N_VSS_Mn8@2197_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2196 N_OUT8_Mn8@2196_d N_OUT7_Mn8@2196_g N_VSS_Mn8@2196_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2197 N_OUT8_Mp8@2197_d N_OUT7_Mp8@2197_g N_VDD_Mp8@2197_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2196 N_OUT8_Mp8@2196_d N_OUT7_Mp8@2196_g N_VDD_Mp8@2196_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2195 N_OUT8_Mn8@2195_d N_OUT7_Mn8@2195_g N_VSS_Mn8@2195_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2194 N_OUT8_Mn8@2194_d N_OUT7_Mn8@2194_g N_VSS_Mn8@2194_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2195 N_OUT8_Mp8@2195_d N_OUT7_Mp8@2195_g N_VDD_Mp8@2195_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2194 N_OUT8_Mp8@2194_d N_OUT7_Mp8@2194_g N_VDD_Mp8@2194_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2193 N_OUT8_Mn8@2193_d N_OUT7_Mn8@2193_g N_VSS_Mn8@2193_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2192 N_OUT8_Mn8@2192_d N_OUT7_Mn8@2192_g N_VSS_Mn8@2192_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2193 N_OUT8_Mp8@2193_d N_OUT7_Mp8@2193_g N_VDD_Mp8@2193_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2192 N_OUT8_Mp8@2192_d N_OUT7_Mp8@2192_g N_VDD_Mp8@2192_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2191 N_OUT8_Mn8@2191_d N_OUT7_Mn8@2191_g N_VSS_Mn8@2191_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2190 N_OUT8_Mn8@2190_d N_OUT7_Mn8@2190_g N_VSS_Mn8@2190_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2191 N_OUT8_Mp8@2191_d N_OUT7_Mp8@2191_g N_VDD_Mp8@2191_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2190 N_OUT8_Mp8@2190_d N_OUT7_Mp8@2190_g N_VDD_Mp8@2190_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2189 N_OUT8_Mn8@2189_d N_OUT7_Mn8@2189_g N_VSS_Mn8@2189_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2188 N_OUT8_Mn8@2188_d N_OUT7_Mn8@2188_g N_VSS_Mn8@2188_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2189 N_OUT8_Mp8@2189_d N_OUT7_Mp8@2189_g N_VDD_Mp8@2189_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2188 N_OUT8_Mp8@2188_d N_OUT7_Mp8@2188_g N_VDD_Mp8@2188_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2187 N_OUT8_Mn8@2187_d N_OUT7_Mn8@2187_g N_VSS_Mn8@2187_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2186 N_OUT8_Mn8@2186_d N_OUT7_Mn8@2186_g N_VSS_Mn8@2186_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2187 N_OUT8_Mp8@2187_d N_OUT7_Mp8@2187_g N_VDD_Mp8@2187_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2186 N_OUT8_Mp8@2186_d N_OUT7_Mp8@2186_g N_VDD_Mp8@2186_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2185 N_OUT8_Mn8@2185_d N_OUT7_Mn8@2185_g N_VSS_Mn8@2185_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2184 N_OUT8_Mn8@2184_d N_OUT7_Mn8@2184_g N_VSS_Mn8@2184_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2185 N_OUT8_Mp8@2185_d N_OUT7_Mp8@2185_g N_VDD_Mp8@2185_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2184 N_OUT8_Mp8@2184_d N_OUT7_Mp8@2184_g N_VDD_Mp8@2184_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2183 N_OUT8_Mn8@2183_d N_OUT7_Mn8@2183_g N_VSS_Mn8@2183_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2182 N_OUT8_Mn8@2182_d N_OUT7_Mn8@2182_g N_VSS_Mn8@2182_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2183 N_OUT8_Mp8@2183_d N_OUT7_Mp8@2183_g N_VDD_Mp8@2183_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2182 N_OUT8_Mp8@2182_d N_OUT7_Mp8@2182_g N_VDD_Mp8@2182_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2181 N_OUT8_Mn8@2181_d N_OUT7_Mn8@2181_g N_VSS_Mn8@2181_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2180 N_OUT8_Mn8@2180_d N_OUT7_Mn8@2180_g N_VSS_Mn8@2180_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2181 N_OUT8_Mp8@2181_d N_OUT7_Mp8@2181_g N_VDD_Mp8@2181_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2180 N_OUT8_Mp8@2180_d N_OUT7_Mp8@2180_g N_VDD_Mp8@2180_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2179 N_OUT8_Mn8@2179_d N_OUT7_Mn8@2179_g N_VSS_Mn8@2179_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2178 N_OUT8_Mn8@2178_d N_OUT7_Mn8@2178_g N_VSS_Mn8@2178_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2179 N_OUT8_Mp8@2179_d N_OUT7_Mp8@2179_g N_VDD_Mp8@2179_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2178 N_OUT8_Mp8@2178_d N_OUT7_Mp8@2178_g N_VDD_Mp8@2178_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2177 N_OUT8_Mn8@2177_d N_OUT7_Mn8@2177_g N_VSS_Mn8@2177_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2176 N_OUT8_Mn8@2176_d N_OUT7_Mn8@2176_g N_VSS_Mn8@2176_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2177 N_OUT8_Mp8@2177_d N_OUT7_Mp8@2177_g N_VDD_Mp8@2177_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2176 N_OUT8_Mp8@2176_d N_OUT7_Mp8@2176_g N_VDD_Mp8@2176_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2175 N_OUT8_Mn8@2175_d N_OUT7_Mn8@2175_g N_VSS_Mn8@2175_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2174 N_OUT8_Mn8@2174_d N_OUT7_Mn8@2174_g N_VSS_Mn8@2174_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2175 N_OUT8_Mp8@2175_d N_OUT7_Mp8@2175_g N_VDD_Mp8@2175_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2174 N_OUT8_Mp8@2174_d N_OUT7_Mp8@2174_g N_VDD_Mp8@2174_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2173 N_OUT8_Mn8@2173_d N_OUT7_Mn8@2173_g N_VSS_Mn8@2173_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2172 N_OUT8_Mn8@2172_d N_OUT7_Mn8@2172_g N_VSS_Mn8@2172_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2173 N_OUT8_Mp8@2173_d N_OUT7_Mp8@2173_g N_VDD_Mp8@2173_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2172 N_OUT8_Mp8@2172_d N_OUT7_Mp8@2172_g N_VDD_Mp8@2172_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2171 N_OUT8_Mn8@2171_d N_OUT7_Mn8@2171_g N_VSS_Mn8@2171_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2170 N_OUT8_Mn8@2170_d N_OUT7_Mn8@2170_g N_VSS_Mn8@2170_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2171 N_OUT8_Mp8@2171_d N_OUT7_Mp8@2171_g N_VDD_Mp8@2171_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2170 N_OUT8_Mp8@2170_d N_OUT7_Mp8@2170_g N_VDD_Mp8@2170_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2169 N_OUT8_Mn8@2169_d N_OUT7_Mn8@2169_g N_VSS_Mn8@2169_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2168 N_OUT8_Mn8@2168_d N_OUT7_Mn8@2168_g N_VSS_Mn8@2168_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2169 N_OUT8_Mp8@2169_d N_OUT7_Mp8@2169_g N_VDD_Mp8@2169_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2168 N_OUT8_Mp8@2168_d N_OUT7_Mp8@2168_g N_VDD_Mp8@2168_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2167 N_OUT8_Mn8@2167_d N_OUT7_Mn8@2167_g N_VSS_Mn8@2167_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2166 N_OUT8_Mn8@2166_d N_OUT7_Mn8@2166_g N_VSS_Mn8@2166_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2167 N_OUT8_Mp8@2167_d N_OUT7_Mp8@2167_g N_VDD_Mp8@2167_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2166 N_OUT8_Mp8@2166_d N_OUT7_Mp8@2166_g N_VDD_Mp8@2166_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2165 N_OUT8_Mn8@2165_d N_OUT7_Mn8@2165_g N_VSS_Mn8@2165_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2164 N_OUT8_Mn8@2164_d N_OUT7_Mn8@2164_g N_VSS_Mn8@2164_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2165 N_OUT8_Mp8@2165_d N_OUT7_Mp8@2165_g N_VDD_Mp8@2165_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2164 N_OUT8_Mp8@2164_d N_OUT7_Mp8@2164_g N_VDD_Mp8@2164_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2163 N_OUT8_Mn8@2163_d N_OUT7_Mn8@2163_g N_VSS_Mn8@2163_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2162 N_OUT8_Mn8@2162_d N_OUT7_Mn8@2162_g N_VSS_Mn8@2162_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2163 N_OUT8_Mp8@2163_d N_OUT7_Mp8@2163_g N_VDD_Mp8@2163_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2162 N_OUT8_Mp8@2162_d N_OUT7_Mp8@2162_g N_VDD_Mp8@2162_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2161 N_OUT8_Mn8@2161_d N_OUT7_Mn8@2161_g N_VSS_Mn8@2161_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2160 N_OUT8_Mn8@2160_d N_OUT7_Mn8@2160_g N_VSS_Mn8@2160_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2161 N_OUT8_Mp8@2161_d N_OUT7_Mp8@2161_g N_VDD_Mp8@2161_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2160 N_OUT8_Mp8@2160_d N_OUT7_Mp8@2160_g N_VDD_Mp8@2160_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2159 N_OUT8_Mn8@2159_d N_OUT7_Mn8@2159_g N_VSS_Mn8@2159_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2158 N_OUT8_Mn8@2158_d N_OUT7_Mn8@2158_g N_VSS_Mn8@2158_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2159 N_OUT8_Mp8@2159_d N_OUT7_Mp8@2159_g N_VDD_Mp8@2159_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2158 N_OUT8_Mp8@2158_d N_OUT7_Mp8@2158_g N_VDD_Mp8@2158_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2157 N_OUT8_Mn8@2157_d N_OUT7_Mn8@2157_g N_VSS_Mn8@2157_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2156 N_OUT8_Mn8@2156_d N_OUT7_Mn8@2156_g N_VSS_Mn8@2156_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2157 N_OUT8_Mp8@2157_d N_OUT7_Mp8@2157_g N_VDD_Mp8@2157_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2156 N_OUT8_Mp8@2156_d N_OUT7_Mp8@2156_g N_VDD_Mp8@2156_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2155 N_OUT8_Mn8@2155_d N_OUT7_Mn8@2155_g N_VSS_Mn8@2155_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2154 N_OUT8_Mn8@2154_d N_OUT7_Mn8@2154_g N_VSS_Mn8@2154_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2155 N_OUT8_Mp8@2155_d N_OUT7_Mp8@2155_g N_VDD_Mp8@2155_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2154 N_OUT8_Mp8@2154_d N_OUT7_Mp8@2154_g N_VDD_Mp8@2154_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2153 N_OUT8_Mn8@2153_d N_OUT7_Mn8@2153_g N_VSS_Mn8@2153_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2152 N_OUT8_Mn8@2152_d N_OUT7_Mn8@2152_g N_VSS_Mn8@2152_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2153 N_OUT8_Mp8@2153_d N_OUT7_Mp8@2153_g N_VDD_Mp8@2153_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2152 N_OUT8_Mp8@2152_d N_OUT7_Mp8@2152_g N_VDD_Mp8@2152_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2151 N_OUT8_Mn8@2151_d N_OUT7_Mn8@2151_g N_VSS_Mn8@2151_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2150 N_OUT8_Mn8@2150_d N_OUT7_Mn8@2150_g N_VSS_Mn8@2150_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2151 N_OUT8_Mp8@2151_d N_OUT7_Mp8@2151_g N_VDD_Mp8@2151_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2150 N_OUT8_Mp8@2150_d N_OUT7_Mp8@2150_g N_VDD_Mp8@2150_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2149 N_OUT8_Mn8@2149_d N_OUT7_Mn8@2149_g N_VSS_Mn8@2149_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2148 N_OUT8_Mn8@2148_d N_OUT7_Mn8@2148_g N_VSS_Mn8@2148_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2149 N_OUT8_Mp8@2149_d N_OUT7_Mp8@2149_g N_VDD_Mp8@2149_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2148 N_OUT8_Mp8@2148_d N_OUT7_Mp8@2148_g N_VDD_Mp8@2148_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2147 N_OUT8_Mn8@2147_d N_OUT7_Mn8@2147_g N_VSS_Mn8@2147_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2146 N_OUT8_Mn8@2146_d N_OUT7_Mn8@2146_g N_VSS_Mn8@2146_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2147 N_OUT8_Mp8@2147_d N_OUT7_Mp8@2147_g N_VDD_Mp8@2147_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2146 N_OUT8_Mp8@2146_d N_OUT7_Mp8@2146_g N_VDD_Mp8@2146_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2145 N_OUT8_Mn8@2145_d N_OUT7_Mn8@2145_g N_VSS_Mn8@2145_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2144 N_OUT8_Mn8@2144_d N_OUT7_Mn8@2144_g N_VSS_Mn8@2144_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2145 N_OUT8_Mp8@2145_d N_OUT7_Mp8@2145_g N_VDD_Mp8@2145_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2144 N_OUT8_Mp8@2144_d N_OUT7_Mp8@2144_g N_VDD_Mp8@2144_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2143 N_OUT8_Mn8@2143_d N_OUT7_Mn8@2143_g N_VSS_Mn8@2143_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2142 N_OUT8_Mn8@2142_d N_OUT7_Mn8@2142_g N_VSS_Mn8@2142_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2143 N_OUT8_Mp8@2143_d N_OUT7_Mp8@2143_g N_VDD_Mp8@2143_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2142 N_OUT8_Mp8@2142_d N_OUT7_Mp8@2142_g N_VDD_Mp8@2142_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2141 N_OUT8_Mn8@2141_d N_OUT7_Mn8@2141_g N_VSS_Mn8@2141_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2140 N_OUT8_Mn8@2140_d N_OUT7_Mn8@2140_g N_VSS_Mn8@2140_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2141 N_OUT8_Mp8@2141_d N_OUT7_Mp8@2141_g N_VDD_Mp8@2141_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2140 N_OUT8_Mp8@2140_d N_OUT7_Mp8@2140_g N_VDD_Mp8@2140_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2139 N_OUT8_Mn8@2139_d N_OUT7_Mn8@2139_g N_VSS_Mn8@2139_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2138 N_OUT8_Mn8@2138_d N_OUT7_Mn8@2138_g N_VSS_Mn8@2138_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2139 N_OUT8_Mp8@2139_d N_OUT7_Mp8@2139_g N_VDD_Mp8@2139_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2138 N_OUT8_Mp8@2138_d N_OUT7_Mp8@2138_g N_VDD_Mp8@2138_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2137 N_OUT8_Mn8@2137_d N_OUT7_Mn8@2137_g N_VSS_Mn8@2137_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2136 N_OUT8_Mn8@2136_d N_OUT7_Mn8@2136_g N_VSS_Mn8@2136_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2137 N_OUT8_Mp8@2137_d N_OUT7_Mp8@2137_g N_VDD_Mp8@2137_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2136 N_OUT8_Mp8@2136_d N_OUT7_Mp8@2136_g N_VDD_Mp8@2136_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2135 N_OUT8_Mn8@2135_d N_OUT7_Mn8@2135_g N_VSS_Mn8@2135_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2134 N_OUT8_Mn8@2134_d N_OUT7_Mn8@2134_g N_VSS_Mn8@2134_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2135 N_OUT8_Mp8@2135_d N_OUT7_Mp8@2135_g N_VDD_Mp8@2135_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2134 N_OUT8_Mp8@2134_d N_OUT7_Mp8@2134_g N_VDD_Mp8@2134_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2133 N_OUT8_Mn8@2133_d N_OUT7_Mn8@2133_g N_VSS_Mn8@2133_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2132 N_OUT8_Mn8@2132_d N_OUT7_Mn8@2132_g N_VSS_Mn8@2132_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2133 N_OUT8_Mp8@2133_d N_OUT7_Mp8@2133_g N_VDD_Mp8@2133_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2132 N_OUT8_Mp8@2132_d N_OUT7_Mp8@2132_g N_VDD_Mp8@2132_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2131 N_OUT8_Mn8@2131_d N_OUT7_Mn8@2131_g N_VSS_Mn8@2131_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2130 N_OUT8_Mn8@2130_d N_OUT7_Mn8@2130_g N_VSS_Mn8@2130_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2131 N_OUT8_Mp8@2131_d N_OUT7_Mp8@2131_g N_VDD_Mp8@2131_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2130 N_OUT8_Mp8@2130_d N_OUT7_Mp8@2130_g N_VDD_Mp8@2130_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2129 N_OUT8_Mn8@2129_d N_OUT7_Mn8@2129_g N_VSS_Mn8@2129_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2128 N_OUT8_Mn8@2128_d N_OUT7_Mn8@2128_g N_VSS_Mn8@2128_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2129 N_OUT8_Mp8@2129_d N_OUT7_Mp8@2129_g N_VDD_Mp8@2129_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2128 N_OUT8_Mp8@2128_d N_OUT7_Mp8@2128_g N_VDD_Mp8@2128_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2127 N_OUT8_Mn8@2127_d N_OUT7_Mn8@2127_g N_VSS_Mn8@2127_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2126 N_OUT8_Mn8@2126_d N_OUT7_Mn8@2126_g N_VSS_Mn8@2126_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2127 N_OUT8_Mp8@2127_d N_OUT7_Mp8@2127_g N_VDD_Mp8@2127_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2126 N_OUT8_Mp8@2126_d N_OUT7_Mp8@2126_g N_VDD_Mp8@2126_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2125 N_OUT8_Mn8@2125_d N_OUT7_Mn8@2125_g N_VSS_Mn8@2125_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2124 N_OUT8_Mn8@2124_d N_OUT7_Mn8@2124_g N_VSS_Mn8@2124_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2125 N_OUT8_Mp8@2125_d N_OUT7_Mp8@2125_g N_VDD_Mp8@2125_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2124 N_OUT8_Mp8@2124_d N_OUT7_Mp8@2124_g N_VDD_Mp8@2124_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2123 N_OUT8_Mn8@2123_d N_OUT7_Mn8@2123_g N_VSS_Mn8@2123_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2122 N_OUT8_Mn8@2122_d N_OUT7_Mn8@2122_g N_VSS_Mn8@2122_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2123 N_OUT8_Mp8@2123_d N_OUT7_Mp8@2123_g N_VDD_Mp8@2123_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2122 N_OUT8_Mp8@2122_d N_OUT7_Mp8@2122_g N_VDD_Mp8@2122_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2121 N_OUT8_Mn8@2121_d N_OUT7_Mn8@2121_g N_VSS_Mn8@2121_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2120 N_OUT8_Mn8@2120_d N_OUT7_Mn8@2120_g N_VSS_Mn8@2120_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2121 N_OUT8_Mp8@2121_d N_OUT7_Mp8@2121_g N_VDD_Mp8@2121_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2120 N_OUT8_Mp8@2120_d N_OUT7_Mp8@2120_g N_VDD_Mp8@2120_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2119 N_OUT8_Mn8@2119_d N_OUT7_Mn8@2119_g N_VSS_Mn8@2119_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2118 N_OUT8_Mn8@2118_d N_OUT7_Mn8@2118_g N_VSS_Mn8@2118_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2119 N_OUT8_Mp8@2119_d N_OUT7_Mp8@2119_g N_VDD_Mp8@2119_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2118 N_OUT8_Mp8@2118_d N_OUT7_Mp8@2118_g N_VDD_Mp8@2118_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2117 N_OUT8_Mn8@2117_d N_OUT7_Mn8@2117_g N_VSS_Mn8@2117_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2116 N_OUT8_Mn8@2116_d N_OUT7_Mn8@2116_g N_VSS_Mn8@2116_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2117 N_OUT8_Mp8@2117_d N_OUT7_Mp8@2117_g N_VDD_Mp8@2117_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2116 N_OUT8_Mp8@2116_d N_OUT7_Mp8@2116_g N_VDD_Mp8@2116_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2115 N_OUT8_Mn8@2115_d N_OUT7_Mn8@2115_g N_VSS_Mn8@2115_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2114 N_OUT8_Mn8@2114_d N_OUT7_Mn8@2114_g N_VSS_Mn8@2114_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2115 N_OUT8_Mp8@2115_d N_OUT7_Mp8@2115_g N_VDD_Mp8@2115_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2114 N_OUT8_Mp8@2114_d N_OUT7_Mp8@2114_g N_VDD_Mp8@2114_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2113 N_OUT8_Mn8@2113_d N_OUT7_Mn8@2113_g N_VSS_Mn8@2113_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2112 N_OUT8_Mn8@2112_d N_OUT7_Mn8@2112_g N_VSS_Mn8@2112_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2113 N_OUT8_Mp8@2113_d N_OUT7_Mp8@2113_g N_VDD_Mp8@2113_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2112 N_OUT8_Mp8@2112_d N_OUT7_Mp8@2112_g N_VDD_Mp8@2112_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2111 N_OUT8_Mn8@2111_d N_OUT7_Mn8@2111_g N_VSS_Mn8@2111_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2110 N_OUT8_Mn8@2110_d N_OUT7_Mn8@2110_g N_VSS_Mn8@2110_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2111 N_OUT8_Mp8@2111_d N_OUT7_Mp8@2111_g N_VDD_Mp8@2111_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2110 N_OUT8_Mp8@2110_d N_OUT7_Mp8@2110_g N_VDD_Mp8@2110_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2109 N_OUT8_Mn8@2109_d N_OUT7_Mn8@2109_g N_VSS_Mn8@2109_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2108 N_OUT8_Mn8@2108_d N_OUT7_Mn8@2108_g N_VSS_Mn8@2108_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2109 N_OUT8_Mp8@2109_d N_OUT7_Mp8@2109_g N_VDD_Mp8@2109_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2108 N_OUT8_Mp8@2108_d N_OUT7_Mp8@2108_g N_VDD_Mp8@2108_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2107 N_OUT8_Mn8@2107_d N_OUT7_Mn8@2107_g N_VSS_Mn8@2107_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2106 N_OUT8_Mn8@2106_d N_OUT7_Mn8@2106_g N_VSS_Mn8@2106_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2107 N_OUT8_Mp8@2107_d N_OUT7_Mp8@2107_g N_VDD_Mp8@2107_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2106 N_OUT8_Mp8@2106_d N_OUT7_Mp8@2106_g N_VDD_Mp8@2106_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2105 N_OUT8_Mn8@2105_d N_OUT7_Mn8@2105_g N_VSS_Mn8@2105_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2104 N_OUT8_Mn8@2104_d N_OUT7_Mn8@2104_g N_VSS_Mn8@2104_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2105 N_OUT8_Mp8@2105_d N_OUT7_Mp8@2105_g N_VDD_Mp8@2105_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2104 N_OUT8_Mp8@2104_d N_OUT7_Mp8@2104_g N_VDD_Mp8@2104_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2103 N_OUT8_Mn8@2103_d N_OUT7_Mn8@2103_g N_VSS_Mn8@2103_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2102 N_OUT8_Mn8@2102_d N_OUT7_Mn8@2102_g N_VSS_Mn8@2102_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2103 N_OUT8_Mp8@2103_d N_OUT7_Mp8@2103_g N_VDD_Mp8@2103_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2102 N_OUT8_Mp8@2102_d N_OUT7_Mp8@2102_g N_VDD_Mp8@2102_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2101 N_OUT8_Mn8@2101_d N_OUT7_Mn8@2101_g N_VSS_Mn8@2101_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2100 N_OUT8_Mn8@2100_d N_OUT7_Mn8@2100_g N_VSS_Mn8@2100_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2101 N_OUT8_Mp8@2101_d N_OUT7_Mp8@2101_g N_VDD_Mp8@2101_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2100 N_OUT8_Mp8@2100_d N_OUT7_Mp8@2100_g N_VDD_Mp8@2100_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2099 N_OUT8_Mn8@2099_d N_OUT7_Mn8@2099_g N_VSS_Mn8@2099_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2098 N_OUT8_Mn8@2098_d N_OUT7_Mn8@2098_g N_VSS_Mn8@2098_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2099 N_OUT8_Mp8@2099_d N_OUT7_Mp8@2099_g N_VDD_Mp8@2099_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2098 N_OUT8_Mp8@2098_d N_OUT7_Mp8@2098_g N_VDD_Mp8@2098_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2097 N_OUT8_Mn8@2097_d N_OUT7_Mn8@2097_g N_VSS_Mn8@2097_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2096 N_OUT8_Mn8@2096_d N_OUT7_Mn8@2096_g N_VSS_Mn8@2096_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2097 N_OUT8_Mp8@2097_d N_OUT7_Mp8@2097_g N_VDD_Mp8@2097_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2096 N_OUT8_Mp8@2096_d N_OUT7_Mp8@2096_g N_VDD_Mp8@2096_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2095 N_OUT8_Mn8@2095_d N_OUT7_Mn8@2095_g N_VSS_Mn8@2095_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2094 N_OUT8_Mn8@2094_d N_OUT7_Mn8@2094_g N_VSS_Mn8@2094_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2095 N_OUT8_Mp8@2095_d N_OUT7_Mp8@2095_g N_VDD_Mp8@2095_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2094 N_OUT8_Mp8@2094_d N_OUT7_Mp8@2094_g N_VDD_Mp8@2094_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2093 N_OUT8_Mn8@2093_d N_OUT7_Mn8@2093_g N_VSS_Mn8@2093_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2092 N_OUT8_Mn8@2092_d N_OUT7_Mn8@2092_g N_VSS_Mn8@2092_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2093 N_OUT8_Mp8@2093_d N_OUT7_Mp8@2093_g N_VDD_Mp8@2093_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2092 N_OUT8_Mp8@2092_d N_OUT7_Mp8@2092_g N_VDD_Mp8@2092_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2091 N_OUT8_Mn8@2091_d N_OUT7_Mn8@2091_g N_VSS_Mn8@2091_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2090 N_OUT8_Mn8@2090_d N_OUT7_Mn8@2090_g N_VSS_Mn8@2090_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2091 N_OUT8_Mp8@2091_d N_OUT7_Mp8@2091_g N_VDD_Mp8@2091_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2090 N_OUT8_Mp8@2090_d N_OUT7_Mp8@2090_g N_VDD_Mp8@2090_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2089 N_OUT8_Mn8@2089_d N_OUT7_Mn8@2089_g N_VSS_Mn8@2089_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2088 N_OUT8_Mn8@2088_d N_OUT7_Mn8@2088_g N_VSS_Mn8@2088_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2089 N_OUT8_Mp8@2089_d N_OUT7_Mp8@2089_g N_VDD_Mp8@2089_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2088 N_OUT8_Mp8@2088_d N_OUT7_Mp8@2088_g N_VDD_Mp8@2088_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2087 N_OUT8_Mn8@2087_d N_OUT7_Mn8@2087_g N_VSS_Mn8@2087_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2086 N_OUT8_Mn8@2086_d N_OUT7_Mn8@2086_g N_VSS_Mn8@2086_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2087 N_OUT8_Mp8@2087_d N_OUT7_Mp8@2087_g N_VDD_Mp8@2087_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2086 N_OUT8_Mp8@2086_d N_OUT7_Mp8@2086_g N_VDD_Mp8@2086_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2085 N_OUT8_Mn8@2085_d N_OUT7_Mn8@2085_g N_VSS_Mn8@2085_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2084 N_OUT8_Mn8@2084_d N_OUT7_Mn8@2084_g N_VSS_Mn8@2084_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2085 N_OUT8_Mp8@2085_d N_OUT7_Mp8@2085_g N_VDD_Mp8@2085_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2084 N_OUT8_Mp8@2084_d N_OUT7_Mp8@2084_g N_VDD_Mp8@2084_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2083 N_OUT8_Mn8@2083_d N_OUT7_Mn8@2083_g N_VSS_Mn8@2083_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2082 N_OUT8_Mn8@2082_d N_OUT7_Mn8@2082_g N_VSS_Mn8@2082_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2083 N_OUT8_Mp8@2083_d N_OUT7_Mp8@2083_g N_VDD_Mp8@2083_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2082 N_OUT8_Mp8@2082_d N_OUT7_Mp8@2082_g N_VDD_Mp8@2082_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2081 N_OUT8_Mn8@2081_d N_OUT7_Mn8@2081_g N_VSS_Mn8@2081_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2080 N_OUT8_Mn8@2080_d N_OUT7_Mn8@2080_g N_VSS_Mn8@2080_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2081 N_OUT8_Mp8@2081_d N_OUT7_Mp8@2081_g N_VDD_Mp8@2081_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2080 N_OUT8_Mp8@2080_d N_OUT7_Mp8@2080_g N_VDD_Mp8@2080_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2079 N_OUT8_Mn8@2079_d N_OUT7_Mn8@2079_g N_VSS_Mn8@2079_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2078 N_OUT8_Mn8@2078_d N_OUT7_Mn8@2078_g N_VSS_Mn8@2078_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2079 N_OUT8_Mp8@2079_d N_OUT7_Mp8@2079_g N_VDD_Mp8@2079_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2078 N_OUT8_Mp8@2078_d N_OUT7_Mp8@2078_g N_VDD_Mp8@2078_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2077 N_OUT8_Mn8@2077_d N_OUT7_Mn8@2077_g N_VSS_Mn8@2077_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2076 N_OUT8_Mn8@2076_d N_OUT7_Mn8@2076_g N_VSS_Mn8@2076_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2077 N_OUT8_Mp8@2077_d N_OUT7_Mp8@2077_g N_VDD_Mp8@2077_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2076 N_OUT8_Mp8@2076_d N_OUT7_Mp8@2076_g N_VDD_Mp8@2076_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2075 N_OUT8_Mn8@2075_d N_OUT7_Mn8@2075_g N_VSS_Mn8@2075_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2074 N_OUT8_Mn8@2074_d N_OUT7_Mn8@2074_g N_VSS_Mn8@2074_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2075 N_OUT8_Mp8@2075_d N_OUT7_Mp8@2075_g N_VDD_Mp8@2075_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2074 N_OUT8_Mp8@2074_d N_OUT7_Mp8@2074_g N_VDD_Mp8@2074_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2073 N_OUT8_Mn8@2073_d N_OUT7_Mn8@2073_g N_VSS_Mn8@2073_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2072 N_OUT8_Mn8@2072_d N_OUT7_Mn8@2072_g N_VSS_Mn8@2072_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2073 N_OUT8_Mp8@2073_d N_OUT7_Mp8@2073_g N_VDD_Mp8@2073_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2072 N_OUT8_Mp8@2072_d N_OUT7_Mp8@2072_g N_VDD_Mp8@2072_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2071 N_OUT8_Mn8@2071_d N_OUT7_Mn8@2071_g N_VSS_Mn8@2071_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2070 N_OUT8_Mn8@2070_d N_OUT7_Mn8@2070_g N_VSS_Mn8@2070_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2071 N_OUT8_Mp8@2071_d N_OUT7_Mp8@2071_g N_VDD_Mp8@2071_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2070 N_OUT8_Mp8@2070_d N_OUT7_Mp8@2070_g N_VDD_Mp8@2070_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2069 N_OUT8_Mn8@2069_d N_OUT7_Mn8@2069_g N_VSS_Mn8@2069_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2068 N_OUT8_Mn8@2068_d N_OUT7_Mn8@2068_g N_VSS_Mn8@2068_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2069 N_OUT8_Mp8@2069_d N_OUT7_Mp8@2069_g N_VDD_Mp8@2069_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2068 N_OUT8_Mp8@2068_d N_OUT7_Mp8@2068_g N_VDD_Mp8@2068_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2067 N_OUT8_Mn8@2067_d N_OUT7_Mn8@2067_g N_VSS_Mn8@2067_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2066 N_OUT8_Mn8@2066_d N_OUT7_Mn8@2066_g N_VSS_Mn8@2066_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2067 N_OUT8_Mp8@2067_d N_OUT7_Mp8@2067_g N_VDD_Mp8@2067_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2066 N_OUT8_Mp8@2066_d N_OUT7_Mp8@2066_g N_VDD_Mp8@2066_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2065 N_OUT8_Mn8@2065_d N_OUT7_Mn8@2065_g N_VSS_Mn8@2065_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2064 N_OUT8_Mn8@2064_d N_OUT7_Mn8@2064_g N_VSS_Mn8@2064_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2065 N_OUT8_Mp8@2065_d N_OUT7_Mp8@2065_g N_VDD_Mp8@2065_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2064 N_OUT8_Mp8@2064_d N_OUT7_Mp8@2064_g N_VDD_Mp8@2064_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2063 N_OUT8_Mn8@2063_d N_OUT7_Mn8@2063_g N_VSS_Mn8@2063_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2062 N_OUT8_Mn8@2062_d N_OUT7_Mn8@2062_g N_VSS_Mn8@2062_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2063 N_OUT8_Mp8@2063_d N_OUT7_Mp8@2063_g N_VDD_Mp8@2063_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2062 N_OUT8_Mp8@2062_d N_OUT7_Mp8@2062_g N_VDD_Mp8@2062_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2061 N_OUT8_Mn8@2061_d N_OUT7_Mn8@2061_g N_VSS_Mn8@2061_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2060 N_OUT8_Mn8@2060_d N_OUT7_Mn8@2060_g N_VSS_Mn8@2060_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2061 N_OUT8_Mp8@2061_d N_OUT7_Mp8@2061_g N_VDD_Mp8@2061_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2060 N_OUT8_Mp8@2060_d N_OUT7_Mp8@2060_g N_VDD_Mp8@2060_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2059 N_OUT8_Mn8@2059_d N_OUT7_Mn8@2059_g N_VSS_Mn8@2059_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2058 N_OUT8_Mn8@2058_d N_OUT7_Mn8@2058_g N_VSS_Mn8@2058_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2059 N_OUT8_Mp8@2059_d N_OUT7_Mp8@2059_g N_VDD_Mp8@2059_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2058 N_OUT8_Mp8@2058_d N_OUT7_Mp8@2058_g N_VDD_Mp8@2058_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2057 N_OUT8_Mn8@2057_d N_OUT7_Mn8@2057_g N_VSS_Mn8@2057_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2056 N_OUT8_Mn8@2056_d N_OUT7_Mn8@2056_g N_VSS_Mn8@2056_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2057 N_OUT8_Mp8@2057_d N_OUT7_Mp8@2057_g N_VDD_Mp8@2057_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2056 N_OUT8_Mp8@2056_d N_OUT7_Mp8@2056_g N_VDD_Mp8@2056_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2055 N_OUT8_Mn8@2055_d N_OUT7_Mn8@2055_g N_VSS_Mn8@2055_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2054 N_OUT8_Mn8@2054_d N_OUT7_Mn8@2054_g N_VSS_Mn8@2054_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2055 N_OUT8_Mp8@2055_d N_OUT7_Mp8@2055_g N_VDD_Mp8@2055_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2054 N_OUT8_Mp8@2054_d N_OUT7_Mp8@2054_g N_VDD_Mp8@2054_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2053 N_OUT8_Mn8@2053_d N_OUT7_Mn8@2053_g N_VSS_Mn8@2053_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2052 N_OUT8_Mn8@2052_d N_OUT7_Mn8@2052_g N_VSS_Mn8@2052_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2053 N_OUT8_Mp8@2053_d N_OUT7_Mp8@2053_g N_VDD_Mp8@2053_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2052 N_OUT8_Mp8@2052_d N_OUT7_Mp8@2052_g N_VDD_Mp8@2052_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2051 N_OUT8_Mn8@2051_d N_OUT7_Mn8@2051_g N_VSS_Mn8@2051_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2050 N_OUT8_Mn8@2050_d N_OUT7_Mn8@2050_g N_VSS_Mn8@2050_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2051 N_OUT8_Mp8@2051_d N_OUT7_Mp8@2051_g N_VDD_Mp8@2051_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2050 N_OUT8_Mp8@2050_d N_OUT7_Mp8@2050_g N_VDD_Mp8@2050_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2049 N_OUT8_Mn8@2049_d N_OUT7_Mn8@2049_g N_VSS_Mn8@2049_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2048 N_OUT8_Mn8@2048_d N_OUT7_Mn8@2048_g N_VSS_Mn8@2048_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2049 N_OUT8_Mp8@2049_d N_OUT7_Mp8@2049_g N_VDD_Mp8@2049_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2048 N_OUT8_Mp8@2048_d N_OUT7_Mp8@2048_g N_VDD_Mp8@2048_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2047 N_OUT8_Mn8@2047_d N_OUT7_Mn8@2047_g N_VSS_Mn8@2047_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2046 N_OUT8_Mn8@2046_d N_OUT7_Mn8@2046_g N_VSS_Mn8@2046_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2047 N_OUT8_Mp8@2047_d N_OUT7_Mp8@2047_g N_VDD_Mp8@2047_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2046 N_OUT8_Mp8@2046_d N_OUT7_Mp8@2046_g N_VDD_Mp8@2046_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2045 N_OUT8_Mn8@2045_d N_OUT7_Mn8@2045_g N_VSS_Mn8@2045_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2044 N_OUT8_Mn8@2044_d N_OUT7_Mn8@2044_g N_VSS_Mn8@2044_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2045 N_OUT8_Mp8@2045_d N_OUT7_Mp8@2045_g N_VDD_Mp8@2045_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2044 N_OUT8_Mp8@2044_d N_OUT7_Mp8@2044_g N_VDD_Mp8@2044_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2043 N_OUT8_Mn8@2043_d N_OUT7_Mn8@2043_g N_VSS_Mn8@2043_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2042 N_OUT8_Mn8@2042_d N_OUT7_Mn8@2042_g N_VSS_Mn8@2042_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2043 N_OUT8_Mp8@2043_d N_OUT7_Mp8@2043_g N_VDD_Mp8@2043_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2042 N_OUT8_Mp8@2042_d N_OUT7_Mp8@2042_g N_VDD_Mp8@2042_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2041 N_OUT8_Mn8@2041_d N_OUT7_Mn8@2041_g N_VSS_Mn8@2041_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2040 N_OUT8_Mn8@2040_d N_OUT7_Mn8@2040_g N_VSS_Mn8@2040_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2041 N_OUT8_Mp8@2041_d N_OUT7_Mp8@2041_g N_VDD_Mp8@2041_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2040 N_OUT8_Mp8@2040_d N_OUT7_Mp8@2040_g N_VDD_Mp8@2040_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2039 N_OUT8_Mn8@2039_d N_OUT7_Mn8@2039_g N_VSS_Mn8@2039_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2038 N_OUT8_Mn8@2038_d N_OUT7_Mn8@2038_g N_VSS_Mn8@2038_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2039 N_OUT8_Mp8@2039_d N_OUT7_Mp8@2039_g N_VDD_Mp8@2039_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2038 N_OUT8_Mp8@2038_d N_OUT7_Mp8@2038_g N_VDD_Mp8@2038_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2037 N_OUT8_Mn8@2037_d N_OUT7_Mn8@2037_g N_VSS_Mn8@2037_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2036 N_OUT8_Mn8@2036_d N_OUT7_Mn8@2036_g N_VSS_Mn8@2036_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2037 N_OUT8_Mp8@2037_d N_OUT7_Mp8@2037_g N_VDD_Mp8@2037_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2036 N_OUT8_Mp8@2036_d N_OUT7_Mp8@2036_g N_VDD_Mp8@2036_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2035 N_OUT8_Mn8@2035_d N_OUT7_Mn8@2035_g N_VSS_Mn8@2035_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2034 N_OUT8_Mn8@2034_d N_OUT7_Mn8@2034_g N_VSS_Mn8@2034_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2035 N_OUT8_Mp8@2035_d N_OUT7_Mp8@2035_g N_VDD_Mp8@2035_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2034 N_OUT8_Mp8@2034_d N_OUT7_Mp8@2034_g N_VDD_Mp8@2034_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2033 N_OUT8_Mn8@2033_d N_OUT7_Mn8@2033_g N_VSS_Mn8@2033_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2032 N_OUT8_Mn8@2032_d N_OUT7_Mn8@2032_g N_VSS_Mn8@2032_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2033 N_OUT8_Mp8@2033_d N_OUT7_Mp8@2033_g N_VDD_Mp8@2033_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2032 N_OUT8_Mp8@2032_d N_OUT7_Mp8@2032_g N_VDD_Mp8@2032_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2031 N_OUT8_Mn8@2031_d N_OUT7_Mn8@2031_g N_VSS_Mn8@2031_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2030 N_OUT8_Mn8@2030_d N_OUT7_Mn8@2030_g N_VSS_Mn8@2030_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2031 N_OUT8_Mp8@2031_d N_OUT7_Mp8@2031_g N_VDD_Mp8@2031_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2030 N_OUT8_Mp8@2030_d N_OUT7_Mp8@2030_g N_VDD_Mp8@2030_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2029 N_OUT8_Mn8@2029_d N_OUT7_Mn8@2029_g N_VSS_Mn8@2029_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2028 N_OUT8_Mn8@2028_d N_OUT7_Mn8@2028_g N_VSS_Mn8@2028_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2029 N_OUT8_Mp8@2029_d N_OUT7_Mp8@2029_g N_VDD_Mp8@2029_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2028 N_OUT8_Mp8@2028_d N_OUT7_Mp8@2028_g N_VDD_Mp8@2028_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2027 N_OUT8_Mn8@2027_d N_OUT7_Mn8@2027_g N_VSS_Mn8@2027_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2026 N_OUT8_Mn8@2026_d N_OUT7_Mn8@2026_g N_VSS_Mn8@2026_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2027 N_OUT8_Mp8@2027_d N_OUT7_Mp8@2027_g N_VDD_Mp8@2027_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2026 N_OUT8_Mp8@2026_d N_OUT7_Mp8@2026_g N_VDD_Mp8@2026_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2025 N_OUT8_Mn8@2025_d N_OUT7_Mn8@2025_g N_VSS_Mn8@2025_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2024 N_OUT8_Mn8@2024_d N_OUT7_Mn8@2024_g N_VSS_Mn8@2024_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2025 N_OUT8_Mp8@2025_d N_OUT7_Mp8@2025_g N_VDD_Mp8@2025_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2024 N_OUT8_Mp8@2024_d N_OUT7_Mp8@2024_g N_VDD_Mp8@2024_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2023 N_OUT8_Mn8@2023_d N_OUT7_Mn8@2023_g N_VSS_Mn8@2023_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2022 N_OUT8_Mn8@2022_d N_OUT7_Mn8@2022_g N_VSS_Mn8@2022_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2023 N_OUT8_Mp8@2023_d N_OUT7_Mp8@2023_g N_VDD_Mp8@2023_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2022 N_OUT8_Mp8@2022_d N_OUT7_Mp8@2022_g N_VDD_Mp8@2022_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2021 N_OUT8_Mn8@2021_d N_OUT7_Mn8@2021_g N_VSS_Mn8@2021_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2020 N_OUT8_Mn8@2020_d N_OUT7_Mn8@2020_g N_VSS_Mn8@2020_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2021 N_OUT8_Mp8@2021_d N_OUT7_Mp8@2021_g N_VDD_Mp8@2021_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2020 N_OUT8_Mp8@2020_d N_OUT7_Mp8@2020_g N_VDD_Mp8@2020_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2019 N_OUT8_Mn8@2019_d N_OUT7_Mn8@2019_g N_VSS_Mn8@2019_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2018 N_OUT8_Mn8@2018_d N_OUT7_Mn8@2018_g N_VSS_Mn8@2018_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2019 N_OUT8_Mp8@2019_d N_OUT7_Mp8@2019_g N_VDD_Mp8@2019_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2018 N_OUT8_Mp8@2018_d N_OUT7_Mp8@2018_g N_VDD_Mp8@2018_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2017 N_OUT8_Mn8@2017_d N_OUT7_Mn8@2017_g N_VSS_Mn8@2017_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2016 N_OUT8_Mn8@2016_d N_OUT7_Mn8@2016_g N_VSS_Mn8@2016_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2017 N_OUT8_Mp8@2017_d N_OUT7_Mp8@2017_g N_VDD_Mp8@2017_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2016 N_OUT8_Mp8@2016_d N_OUT7_Mp8@2016_g N_VDD_Mp8@2016_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2015 N_OUT8_Mn8@2015_d N_OUT7_Mn8@2015_g N_VSS_Mn8@2015_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2014 N_OUT8_Mn8@2014_d N_OUT7_Mn8@2014_g N_VSS_Mn8@2014_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2015 N_OUT8_Mp8@2015_d N_OUT7_Mp8@2015_g N_VDD_Mp8@2015_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2014 N_OUT8_Mp8@2014_d N_OUT7_Mp8@2014_g N_VDD_Mp8@2014_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2013 N_OUT8_Mn8@2013_d N_OUT7_Mn8@2013_g N_VSS_Mn8@2013_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2012 N_OUT8_Mn8@2012_d N_OUT7_Mn8@2012_g N_VSS_Mn8@2012_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2013 N_OUT8_Mp8@2013_d N_OUT7_Mp8@2013_g N_VDD_Mp8@2013_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2012 N_OUT8_Mp8@2012_d N_OUT7_Mp8@2012_g N_VDD_Mp8@2012_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2011 N_OUT8_Mn8@2011_d N_OUT7_Mn8@2011_g N_VSS_Mn8@2011_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2010 N_OUT8_Mn8@2010_d N_OUT7_Mn8@2010_g N_VSS_Mn8@2010_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2011 N_OUT8_Mp8@2011_d N_OUT7_Mp8@2011_g N_VDD_Mp8@2011_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2010 N_OUT8_Mp8@2010_d N_OUT7_Mp8@2010_g N_VDD_Mp8@2010_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2009 N_OUT8_Mn8@2009_d N_OUT7_Mn8@2009_g N_VSS_Mn8@2009_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2008 N_OUT8_Mn8@2008_d N_OUT7_Mn8@2008_g N_VSS_Mn8@2008_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2009 N_OUT8_Mp8@2009_d N_OUT7_Mp8@2009_g N_VDD_Mp8@2009_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2008 N_OUT8_Mp8@2008_d N_OUT7_Mp8@2008_g N_VDD_Mp8@2008_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2007 N_OUT8_Mn8@2007_d N_OUT7_Mn8@2007_g N_VSS_Mn8@2007_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2006 N_OUT8_Mn8@2006_d N_OUT7_Mn8@2006_g N_VSS_Mn8@2006_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2007 N_OUT8_Mp8@2007_d N_OUT7_Mp8@2007_g N_VDD_Mp8@2007_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2006 N_OUT8_Mp8@2006_d N_OUT7_Mp8@2006_g N_VDD_Mp8@2006_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2005 N_OUT8_Mn8@2005_d N_OUT7_Mn8@2005_g N_VSS_Mn8@2005_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2004 N_OUT8_Mn8@2004_d N_OUT7_Mn8@2004_g N_VSS_Mn8@2004_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2005 N_OUT8_Mp8@2005_d N_OUT7_Mp8@2005_g N_VDD_Mp8@2005_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2004 N_OUT8_Mp8@2004_d N_OUT7_Mp8@2004_g N_VDD_Mp8@2004_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2003 N_OUT8_Mn8@2003_d N_OUT7_Mn8@2003_g N_VSS_Mn8@2003_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2002 N_OUT8_Mn8@2002_d N_OUT7_Mn8@2002_g N_VSS_Mn8@2002_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2003 N_OUT8_Mp8@2003_d N_OUT7_Mp8@2003_g N_VDD_Mp8@2003_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2002 N_OUT8_Mp8@2002_d N_OUT7_Mp8@2002_g N_VDD_Mp8@2002_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@2001 N_OUT8_Mn8@2001_d N_OUT7_Mn8@2001_g N_VSS_Mn8@2001_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2000 N_OUT8_Mn8@2000_d N_OUT7_Mn8@2000_g N_VSS_Mn8@2000_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@2001 N_OUT8_Mp8@2001_d N_OUT7_Mp8@2001_g N_VDD_Mp8@2001_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2000 N_OUT8_Mp8@2000_d N_OUT7_Mp8@2000_g N_VDD_Mp8@2000_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1999 N_OUT8_Mn8@1999_d N_OUT7_Mn8@1999_g N_VSS_Mn8@1999_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1998 N_OUT8_Mn8@1998_d N_OUT7_Mn8@1998_g N_VSS_Mn8@1998_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1999 N_OUT8_Mp8@1999_d N_OUT7_Mp8@1999_g N_VDD_Mp8@1999_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1998 N_OUT8_Mp8@1998_d N_OUT7_Mp8@1998_g N_VDD_Mp8@1998_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1997 N_OUT8_Mn8@1997_d N_OUT7_Mn8@1997_g N_VSS_Mn8@1997_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1996 N_OUT8_Mn8@1996_d N_OUT7_Mn8@1996_g N_VSS_Mn8@1996_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1997 N_OUT8_Mp8@1997_d N_OUT7_Mp8@1997_g N_VDD_Mp8@1997_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1996 N_OUT8_Mp8@1996_d N_OUT7_Mp8@1996_g N_VDD_Mp8@1996_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1995 N_OUT8_Mn8@1995_d N_OUT7_Mn8@1995_g N_VSS_Mn8@1995_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1994 N_OUT8_Mn8@1994_d N_OUT7_Mn8@1994_g N_VSS_Mn8@1994_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1995 N_OUT8_Mp8@1995_d N_OUT7_Mp8@1995_g N_VDD_Mp8@1995_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1994 N_OUT8_Mp8@1994_d N_OUT7_Mp8@1994_g N_VDD_Mp8@1994_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1993 N_OUT8_Mn8@1993_d N_OUT7_Mn8@1993_g N_VSS_Mn8@1993_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1992 N_OUT8_Mn8@1992_d N_OUT7_Mn8@1992_g N_VSS_Mn8@1992_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1993 N_OUT8_Mp8@1993_d N_OUT7_Mp8@1993_g N_VDD_Mp8@1993_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1992 N_OUT8_Mp8@1992_d N_OUT7_Mp8@1992_g N_VDD_Mp8@1992_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1991 N_OUT8_Mn8@1991_d N_OUT7_Mn8@1991_g N_VSS_Mn8@1991_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1990 N_OUT8_Mn8@1990_d N_OUT7_Mn8@1990_g N_VSS_Mn8@1990_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1991 N_OUT8_Mp8@1991_d N_OUT7_Mp8@1991_g N_VDD_Mp8@1991_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1990 N_OUT8_Mp8@1990_d N_OUT7_Mp8@1990_g N_VDD_Mp8@1990_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1989 N_OUT8_Mn8@1989_d N_OUT7_Mn8@1989_g N_VSS_Mn8@1989_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1988 N_OUT8_Mn8@1988_d N_OUT7_Mn8@1988_g N_VSS_Mn8@1988_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1989 N_OUT8_Mp8@1989_d N_OUT7_Mp8@1989_g N_VDD_Mp8@1989_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1988 N_OUT8_Mp8@1988_d N_OUT7_Mp8@1988_g N_VDD_Mp8@1988_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1987 N_OUT8_Mn8@1987_d N_OUT7_Mn8@1987_g N_VSS_Mn8@1987_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1986 N_OUT8_Mn8@1986_d N_OUT7_Mn8@1986_g N_VSS_Mn8@1986_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1987 N_OUT8_Mp8@1987_d N_OUT7_Mp8@1987_g N_VDD_Mp8@1987_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1986 N_OUT8_Mp8@1986_d N_OUT7_Mp8@1986_g N_VDD_Mp8@1986_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1985 N_OUT8_Mn8@1985_d N_OUT7_Mn8@1985_g N_VSS_Mn8@1985_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1984 N_OUT8_Mn8@1984_d N_OUT7_Mn8@1984_g N_VSS_Mn8@1984_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1985 N_OUT8_Mp8@1985_d N_OUT7_Mp8@1985_g N_VDD_Mp8@1985_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1984 N_OUT8_Mp8@1984_d N_OUT7_Mp8@1984_g N_VDD_Mp8@1984_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1983 N_OUT8_Mn8@1983_d N_OUT7_Mn8@1983_g N_VSS_Mn8@1983_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1982 N_OUT8_Mn8@1982_d N_OUT7_Mn8@1982_g N_VSS_Mn8@1982_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1983 N_OUT8_Mp8@1983_d N_OUT7_Mp8@1983_g N_VDD_Mp8@1983_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1982 N_OUT8_Mp8@1982_d N_OUT7_Mp8@1982_g N_VDD_Mp8@1982_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1981 N_OUT8_Mn8@1981_d N_OUT7_Mn8@1981_g N_VSS_Mn8@1981_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1980 N_OUT8_Mn8@1980_d N_OUT7_Mn8@1980_g N_VSS_Mn8@1980_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1981 N_OUT8_Mp8@1981_d N_OUT7_Mp8@1981_g N_VDD_Mp8@1981_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1980 N_OUT8_Mp8@1980_d N_OUT7_Mp8@1980_g N_VDD_Mp8@1980_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1979 N_OUT8_Mn8@1979_d N_OUT7_Mn8@1979_g N_VSS_Mn8@1979_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1978 N_OUT8_Mn8@1978_d N_OUT7_Mn8@1978_g N_VSS_Mn8@1978_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1979 N_OUT8_Mp8@1979_d N_OUT7_Mp8@1979_g N_VDD_Mp8@1979_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1978 N_OUT8_Mp8@1978_d N_OUT7_Mp8@1978_g N_VDD_Mp8@1978_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1977 N_OUT8_Mn8@1977_d N_OUT7_Mn8@1977_g N_VSS_Mn8@1977_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1976 N_OUT8_Mn8@1976_d N_OUT7_Mn8@1976_g N_VSS_Mn8@1976_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1977 N_OUT8_Mp8@1977_d N_OUT7_Mp8@1977_g N_VDD_Mp8@1977_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1976 N_OUT8_Mp8@1976_d N_OUT7_Mp8@1976_g N_VDD_Mp8@1976_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1975 N_OUT8_Mn8@1975_d N_OUT7_Mn8@1975_g N_VSS_Mn8@1975_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1974 N_OUT8_Mn8@1974_d N_OUT7_Mn8@1974_g N_VSS_Mn8@1974_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1975 N_OUT8_Mp8@1975_d N_OUT7_Mp8@1975_g N_VDD_Mp8@1975_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1974 N_OUT8_Mp8@1974_d N_OUT7_Mp8@1974_g N_VDD_Mp8@1974_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1973 N_OUT8_Mn8@1973_d N_OUT7_Mn8@1973_g N_VSS_Mn8@1973_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1972 N_OUT8_Mn8@1972_d N_OUT7_Mn8@1972_g N_VSS_Mn8@1972_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1973 N_OUT8_Mp8@1973_d N_OUT7_Mp8@1973_g N_VDD_Mp8@1973_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1972 N_OUT8_Mp8@1972_d N_OUT7_Mp8@1972_g N_VDD_Mp8@1972_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1971 N_OUT8_Mn8@1971_d N_OUT7_Mn8@1971_g N_VSS_Mn8@1971_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1970 N_OUT8_Mn8@1970_d N_OUT7_Mn8@1970_g N_VSS_Mn8@1970_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1971 N_OUT8_Mp8@1971_d N_OUT7_Mp8@1971_g N_VDD_Mp8@1971_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1970 N_OUT8_Mp8@1970_d N_OUT7_Mp8@1970_g N_VDD_Mp8@1970_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1969 N_OUT8_Mn8@1969_d N_OUT7_Mn8@1969_g N_VSS_Mn8@1969_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1968 N_OUT8_Mn8@1968_d N_OUT7_Mn8@1968_g N_VSS_Mn8@1968_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1969 N_OUT8_Mp8@1969_d N_OUT7_Mp8@1969_g N_VDD_Mp8@1969_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1968 N_OUT8_Mp8@1968_d N_OUT7_Mp8@1968_g N_VDD_Mp8@1968_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1967 N_OUT8_Mn8@1967_d N_OUT7_Mn8@1967_g N_VSS_Mn8@1967_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1966 N_OUT8_Mn8@1966_d N_OUT7_Mn8@1966_g N_VSS_Mn8@1966_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1967 N_OUT8_Mp8@1967_d N_OUT7_Mp8@1967_g N_VDD_Mp8@1967_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1966 N_OUT8_Mp8@1966_d N_OUT7_Mp8@1966_g N_VDD_Mp8@1966_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1965 N_OUT8_Mn8@1965_d N_OUT7_Mn8@1965_g N_VSS_Mn8@1965_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1964 N_OUT8_Mn8@1964_d N_OUT7_Mn8@1964_g N_VSS_Mn8@1964_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1965 N_OUT8_Mp8@1965_d N_OUT7_Mp8@1965_g N_VDD_Mp8@1965_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1964 N_OUT8_Mp8@1964_d N_OUT7_Mp8@1964_g N_VDD_Mp8@1964_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1963 N_OUT8_Mn8@1963_d N_OUT7_Mn8@1963_g N_VSS_Mn8@1963_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1962 N_OUT8_Mn8@1962_d N_OUT7_Mn8@1962_g N_VSS_Mn8@1962_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1963 N_OUT8_Mp8@1963_d N_OUT7_Mp8@1963_g N_VDD_Mp8@1963_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1962 N_OUT8_Mp8@1962_d N_OUT7_Mp8@1962_g N_VDD_Mp8@1962_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1961 N_OUT8_Mn8@1961_d N_OUT7_Mn8@1961_g N_VSS_Mn8@1961_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1960 N_OUT8_Mn8@1960_d N_OUT7_Mn8@1960_g N_VSS_Mn8@1960_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1961 N_OUT8_Mp8@1961_d N_OUT7_Mp8@1961_g N_VDD_Mp8@1961_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1960 N_OUT8_Mp8@1960_d N_OUT7_Mp8@1960_g N_VDD_Mp8@1960_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1959 N_OUT8_Mn8@1959_d N_OUT7_Mn8@1959_g N_VSS_Mn8@1959_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1958 N_OUT8_Mn8@1958_d N_OUT7_Mn8@1958_g N_VSS_Mn8@1958_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1959 N_OUT8_Mp8@1959_d N_OUT7_Mp8@1959_g N_VDD_Mp8@1959_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1958 N_OUT8_Mp8@1958_d N_OUT7_Mp8@1958_g N_VDD_Mp8@1958_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1957 N_OUT8_Mn8@1957_d N_OUT7_Mn8@1957_g N_VSS_Mn8@1957_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1956 N_OUT8_Mn8@1956_d N_OUT7_Mn8@1956_g N_VSS_Mn8@1956_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1957 N_OUT8_Mp8@1957_d N_OUT7_Mp8@1957_g N_VDD_Mp8@1957_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1956 N_OUT8_Mp8@1956_d N_OUT7_Mp8@1956_g N_VDD_Mp8@1956_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1955 N_OUT8_Mn8@1955_d N_OUT7_Mn8@1955_g N_VSS_Mn8@1955_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1954 N_OUT8_Mn8@1954_d N_OUT7_Mn8@1954_g N_VSS_Mn8@1954_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1955 N_OUT8_Mp8@1955_d N_OUT7_Mp8@1955_g N_VDD_Mp8@1955_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1954 N_OUT8_Mp8@1954_d N_OUT7_Mp8@1954_g N_VDD_Mp8@1954_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1953 N_OUT8_Mn8@1953_d N_OUT7_Mn8@1953_g N_VSS_Mn8@1953_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1952 N_OUT8_Mn8@1952_d N_OUT7_Mn8@1952_g N_VSS_Mn8@1952_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1953 N_OUT8_Mp8@1953_d N_OUT7_Mp8@1953_g N_VDD_Mp8@1953_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1952 N_OUT8_Mp8@1952_d N_OUT7_Mp8@1952_g N_VDD_Mp8@1952_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1951 N_OUT8_Mn8@1951_d N_OUT7_Mn8@1951_g N_VSS_Mn8@1951_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1950 N_OUT8_Mn8@1950_d N_OUT7_Mn8@1950_g N_VSS_Mn8@1950_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1951 N_OUT8_Mp8@1951_d N_OUT7_Mp8@1951_g N_VDD_Mp8@1951_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1950 N_OUT8_Mp8@1950_d N_OUT7_Mp8@1950_g N_VDD_Mp8@1950_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1949 N_OUT8_Mn8@1949_d N_OUT7_Mn8@1949_g N_VSS_Mn8@1949_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1948 N_OUT8_Mn8@1948_d N_OUT7_Mn8@1948_g N_VSS_Mn8@1948_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1949 N_OUT8_Mp8@1949_d N_OUT7_Mp8@1949_g N_VDD_Mp8@1949_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1948 N_OUT8_Mp8@1948_d N_OUT7_Mp8@1948_g N_VDD_Mp8@1948_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1947 N_OUT8_Mn8@1947_d N_OUT7_Mn8@1947_g N_VSS_Mn8@1947_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1946 N_OUT8_Mn8@1946_d N_OUT7_Mn8@1946_g N_VSS_Mn8@1946_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1947 N_OUT8_Mp8@1947_d N_OUT7_Mp8@1947_g N_VDD_Mp8@1947_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1946 N_OUT8_Mp8@1946_d N_OUT7_Mp8@1946_g N_VDD_Mp8@1946_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1945 N_OUT8_Mn8@1945_d N_OUT7_Mn8@1945_g N_VSS_Mn8@1945_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1944 N_OUT8_Mn8@1944_d N_OUT7_Mn8@1944_g N_VSS_Mn8@1944_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1945 N_OUT8_Mp8@1945_d N_OUT7_Mp8@1945_g N_VDD_Mp8@1945_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1944 N_OUT8_Mp8@1944_d N_OUT7_Mp8@1944_g N_VDD_Mp8@1944_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1943 N_OUT8_Mn8@1943_d N_OUT7_Mn8@1943_g N_VSS_Mn8@1943_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1942 N_OUT8_Mn8@1942_d N_OUT7_Mn8@1942_g N_VSS_Mn8@1942_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1943 N_OUT8_Mp8@1943_d N_OUT7_Mp8@1943_g N_VDD_Mp8@1943_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1942 N_OUT8_Mp8@1942_d N_OUT7_Mp8@1942_g N_VDD_Mp8@1942_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1941 N_OUT8_Mn8@1941_d N_OUT7_Mn8@1941_g N_VSS_Mn8@1941_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1940 N_OUT8_Mn8@1940_d N_OUT7_Mn8@1940_g N_VSS_Mn8@1940_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1941 N_OUT8_Mp8@1941_d N_OUT7_Mp8@1941_g N_VDD_Mp8@1941_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1940 N_OUT8_Mp8@1940_d N_OUT7_Mp8@1940_g N_VDD_Mp8@1940_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1939 N_OUT8_Mn8@1939_d N_OUT7_Mn8@1939_g N_VSS_Mn8@1939_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1938 N_OUT8_Mn8@1938_d N_OUT7_Mn8@1938_g N_VSS_Mn8@1938_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1939 N_OUT8_Mp8@1939_d N_OUT7_Mp8@1939_g N_VDD_Mp8@1939_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1938 N_OUT8_Mp8@1938_d N_OUT7_Mp8@1938_g N_VDD_Mp8@1938_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1937 N_OUT8_Mn8@1937_d N_OUT7_Mn8@1937_g N_VSS_Mn8@1937_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1936 N_OUT8_Mn8@1936_d N_OUT7_Mn8@1936_g N_VSS_Mn8@1936_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1937 N_OUT8_Mp8@1937_d N_OUT7_Mp8@1937_g N_VDD_Mp8@1937_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1936 N_OUT8_Mp8@1936_d N_OUT7_Mp8@1936_g N_VDD_Mp8@1936_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1935 N_OUT8_Mn8@1935_d N_OUT7_Mn8@1935_g N_VSS_Mn8@1935_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1934 N_OUT8_Mn8@1934_d N_OUT7_Mn8@1934_g N_VSS_Mn8@1934_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1935 N_OUT8_Mp8@1935_d N_OUT7_Mp8@1935_g N_VDD_Mp8@1935_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1934 N_OUT8_Mp8@1934_d N_OUT7_Mp8@1934_g N_VDD_Mp8@1934_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1933 N_OUT8_Mn8@1933_d N_OUT7_Mn8@1933_g N_VSS_Mn8@1933_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1932 N_OUT8_Mn8@1932_d N_OUT7_Mn8@1932_g N_VSS_Mn8@1932_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1933 N_OUT8_Mp8@1933_d N_OUT7_Mp8@1933_g N_VDD_Mp8@1933_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1932 N_OUT8_Mp8@1932_d N_OUT7_Mp8@1932_g N_VDD_Mp8@1932_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1931 N_OUT8_Mn8@1931_d N_OUT7_Mn8@1931_g N_VSS_Mn8@1931_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1930 N_OUT8_Mn8@1930_d N_OUT7_Mn8@1930_g N_VSS_Mn8@1930_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1931 N_OUT8_Mp8@1931_d N_OUT7_Mp8@1931_g N_VDD_Mp8@1931_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1930 N_OUT8_Mp8@1930_d N_OUT7_Mp8@1930_g N_VDD_Mp8@1930_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1929 N_OUT8_Mn8@1929_d N_OUT7_Mn8@1929_g N_VSS_Mn8@1929_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1928 N_OUT8_Mn8@1928_d N_OUT7_Mn8@1928_g N_VSS_Mn8@1928_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1929 N_OUT8_Mp8@1929_d N_OUT7_Mp8@1929_g N_VDD_Mp8@1929_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1928 N_OUT8_Mp8@1928_d N_OUT7_Mp8@1928_g N_VDD_Mp8@1928_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1927 N_OUT8_Mn8@1927_d N_OUT7_Mn8@1927_g N_VSS_Mn8@1927_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1926 N_OUT8_Mn8@1926_d N_OUT7_Mn8@1926_g N_VSS_Mn8@1926_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1927 N_OUT8_Mp8@1927_d N_OUT7_Mp8@1927_g N_VDD_Mp8@1927_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1926 N_OUT8_Mp8@1926_d N_OUT7_Mp8@1926_g N_VDD_Mp8@1926_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1925 N_OUT8_Mn8@1925_d N_OUT7_Mn8@1925_g N_VSS_Mn8@1925_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1924 N_OUT8_Mn8@1924_d N_OUT7_Mn8@1924_g N_VSS_Mn8@1924_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1925 N_OUT8_Mp8@1925_d N_OUT7_Mp8@1925_g N_VDD_Mp8@1925_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1924 N_OUT8_Mp8@1924_d N_OUT7_Mp8@1924_g N_VDD_Mp8@1924_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1923 N_OUT8_Mn8@1923_d N_OUT7_Mn8@1923_g N_VSS_Mn8@1923_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1922 N_OUT8_Mn8@1922_d N_OUT7_Mn8@1922_g N_VSS_Mn8@1922_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1923 N_OUT8_Mp8@1923_d N_OUT7_Mp8@1923_g N_VDD_Mp8@1923_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1922 N_OUT8_Mp8@1922_d N_OUT7_Mp8@1922_g N_VDD_Mp8@1922_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1921 N_OUT8_Mn8@1921_d N_OUT7_Mn8@1921_g N_VSS_Mn8@1921_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1920 N_OUT8_Mn8@1920_d N_OUT7_Mn8@1920_g N_VSS_Mn8@1920_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1921 N_OUT8_Mp8@1921_d N_OUT7_Mp8@1921_g N_VDD_Mp8@1921_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1920 N_OUT8_Mp8@1920_d N_OUT7_Mp8@1920_g N_VDD_Mp8@1920_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1919 N_OUT8_Mn8@1919_d N_OUT7_Mn8@1919_g N_VSS_Mn8@1919_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1918 N_OUT8_Mn8@1918_d N_OUT7_Mn8@1918_g N_VSS_Mn8@1918_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1919 N_OUT8_Mp8@1919_d N_OUT7_Mp8@1919_g N_VDD_Mp8@1919_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1918 N_OUT8_Mp8@1918_d N_OUT7_Mp8@1918_g N_VDD_Mp8@1918_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1917 N_OUT8_Mn8@1917_d N_OUT7_Mn8@1917_g N_VSS_Mn8@1917_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1916 N_OUT8_Mn8@1916_d N_OUT7_Mn8@1916_g N_VSS_Mn8@1916_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1917 N_OUT8_Mp8@1917_d N_OUT7_Mp8@1917_g N_VDD_Mp8@1917_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1916 N_OUT8_Mp8@1916_d N_OUT7_Mp8@1916_g N_VDD_Mp8@1916_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1915 N_OUT8_Mn8@1915_d N_OUT7_Mn8@1915_g N_VSS_Mn8@1915_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1914 N_OUT8_Mn8@1914_d N_OUT7_Mn8@1914_g N_VSS_Mn8@1914_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1915 N_OUT8_Mp8@1915_d N_OUT7_Mp8@1915_g N_VDD_Mp8@1915_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1914 N_OUT8_Mp8@1914_d N_OUT7_Mp8@1914_g N_VDD_Mp8@1914_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1913 N_OUT8_Mn8@1913_d N_OUT7_Mn8@1913_g N_VSS_Mn8@1913_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1912 N_OUT8_Mn8@1912_d N_OUT7_Mn8@1912_g N_VSS_Mn8@1912_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1913 N_OUT8_Mp8@1913_d N_OUT7_Mp8@1913_g N_VDD_Mp8@1913_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1912 N_OUT8_Mp8@1912_d N_OUT7_Mp8@1912_g N_VDD_Mp8@1912_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1911 N_OUT8_Mn8@1911_d N_OUT7_Mn8@1911_g N_VSS_Mn8@1911_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1910 N_OUT8_Mn8@1910_d N_OUT7_Mn8@1910_g N_VSS_Mn8@1910_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1911 N_OUT8_Mp8@1911_d N_OUT7_Mp8@1911_g N_VDD_Mp8@1911_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1910 N_OUT8_Mp8@1910_d N_OUT7_Mp8@1910_g N_VDD_Mp8@1910_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1909 N_OUT8_Mn8@1909_d N_OUT7_Mn8@1909_g N_VSS_Mn8@1909_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1908 N_OUT8_Mn8@1908_d N_OUT7_Mn8@1908_g N_VSS_Mn8@1908_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1909 N_OUT8_Mp8@1909_d N_OUT7_Mp8@1909_g N_VDD_Mp8@1909_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1908 N_OUT8_Mp8@1908_d N_OUT7_Mp8@1908_g N_VDD_Mp8@1908_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1907 N_OUT8_Mn8@1907_d N_OUT7_Mn8@1907_g N_VSS_Mn8@1907_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1906 N_OUT8_Mn8@1906_d N_OUT7_Mn8@1906_g N_VSS_Mn8@1906_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1907 N_OUT8_Mp8@1907_d N_OUT7_Mp8@1907_g N_VDD_Mp8@1907_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1906 N_OUT8_Mp8@1906_d N_OUT7_Mp8@1906_g N_VDD_Mp8@1906_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1905 N_OUT8_Mn8@1905_d N_OUT7_Mn8@1905_g N_VSS_Mn8@1905_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1904 N_OUT8_Mn8@1904_d N_OUT7_Mn8@1904_g N_VSS_Mn8@1904_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1905 N_OUT8_Mp8@1905_d N_OUT7_Mp8@1905_g N_VDD_Mp8@1905_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1904 N_OUT8_Mp8@1904_d N_OUT7_Mp8@1904_g N_VDD_Mp8@1904_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1903 N_OUT8_Mn8@1903_d N_OUT7_Mn8@1903_g N_VSS_Mn8@1903_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1902 N_OUT8_Mn8@1902_d N_OUT7_Mn8@1902_g N_VSS_Mn8@1902_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1903 N_OUT8_Mp8@1903_d N_OUT7_Mp8@1903_g N_VDD_Mp8@1903_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1902 N_OUT8_Mp8@1902_d N_OUT7_Mp8@1902_g N_VDD_Mp8@1902_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1901 N_OUT8_Mn8@1901_d N_OUT7_Mn8@1901_g N_VSS_Mn8@1901_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1900 N_OUT8_Mn8@1900_d N_OUT7_Mn8@1900_g N_VSS_Mn8@1900_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1901 N_OUT8_Mp8@1901_d N_OUT7_Mp8@1901_g N_VDD_Mp8@1901_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1900 N_OUT8_Mp8@1900_d N_OUT7_Mp8@1900_g N_VDD_Mp8@1900_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1899 N_OUT8_Mn8@1899_d N_OUT7_Mn8@1899_g N_VSS_Mn8@1899_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1898 N_OUT8_Mn8@1898_d N_OUT7_Mn8@1898_g N_VSS_Mn8@1898_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1899 N_OUT8_Mp8@1899_d N_OUT7_Mp8@1899_g N_VDD_Mp8@1899_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1898 N_OUT8_Mp8@1898_d N_OUT7_Mp8@1898_g N_VDD_Mp8@1898_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1897 N_OUT8_Mn8@1897_d N_OUT7_Mn8@1897_g N_VSS_Mn8@1897_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1896 N_OUT8_Mn8@1896_d N_OUT7_Mn8@1896_g N_VSS_Mn8@1896_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1897 N_OUT8_Mp8@1897_d N_OUT7_Mp8@1897_g N_VDD_Mp8@1897_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1896 N_OUT8_Mp8@1896_d N_OUT7_Mp8@1896_g N_VDD_Mp8@1896_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1895 N_OUT8_Mn8@1895_d N_OUT7_Mn8@1895_g N_VSS_Mn8@1895_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1894 N_OUT8_Mn8@1894_d N_OUT7_Mn8@1894_g N_VSS_Mn8@1894_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1895 N_OUT8_Mp8@1895_d N_OUT7_Mp8@1895_g N_VDD_Mp8@1895_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1894 N_OUT8_Mp8@1894_d N_OUT7_Mp8@1894_g N_VDD_Mp8@1894_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1893 N_OUT8_Mn8@1893_d N_OUT7_Mn8@1893_g N_VSS_Mn8@1893_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1892 N_OUT8_Mn8@1892_d N_OUT7_Mn8@1892_g N_VSS_Mn8@1892_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1893 N_OUT8_Mp8@1893_d N_OUT7_Mp8@1893_g N_VDD_Mp8@1893_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1892 N_OUT8_Mp8@1892_d N_OUT7_Mp8@1892_g N_VDD_Mp8@1892_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1891 N_OUT8_Mn8@1891_d N_OUT7_Mn8@1891_g N_VSS_Mn8@1891_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1890 N_OUT8_Mn8@1890_d N_OUT7_Mn8@1890_g N_VSS_Mn8@1890_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1891 N_OUT8_Mp8@1891_d N_OUT7_Mp8@1891_g N_VDD_Mp8@1891_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1890 N_OUT8_Mp8@1890_d N_OUT7_Mp8@1890_g N_VDD_Mp8@1890_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1889 N_OUT8_Mn8@1889_d N_OUT7_Mn8@1889_g N_VSS_Mn8@1889_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1888 N_OUT8_Mn8@1888_d N_OUT7_Mn8@1888_g N_VSS_Mn8@1888_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1889 N_OUT8_Mp8@1889_d N_OUT7_Mp8@1889_g N_VDD_Mp8@1889_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1888 N_OUT8_Mp8@1888_d N_OUT7_Mp8@1888_g N_VDD_Mp8@1888_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1887 N_OUT8_Mn8@1887_d N_OUT7_Mn8@1887_g N_VSS_Mn8@1887_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1886 N_OUT8_Mn8@1886_d N_OUT7_Mn8@1886_g N_VSS_Mn8@1886_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1887 N_OUT8_Mp8@1887_d N_OUT7_Mp8@1887_g N_VDD_Mp8@1887_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1886 N_OUT8_Mp8@1886_d N_OUT7_Mp8@1886_g N_VDD_Mp8@1886_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1885 N_OUT8_Mn8@1885_d N_OUT7_Mn8@1885_g N_VSS_Mn8@1885_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1884 N_OUT8_Mn8@1884_d N_OUT7_Mn8@1884_g N_VSS_Mn8@1884_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1885 N_OUT8_Mp8@1885_d N_OUT7_Mp8@1885_g N_VDD_Mp8@1885_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1884 N_OUT8_Mp8@1884_d N_OUT7_Mp8@1884_g N_VDD_Mp8@1884_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1883 N_OUT8_Mn8@1883_d N_OUT7_Mn8@1883_g N_VSS_Mn8@1883_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1882 N_OUT8_Mn8@1882_d N_OUT7_Mn8@1882_g N_VSS_Mn8@1882_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1883 N_OUT8_Mp8@1883_d N_OUT7_Mp8@1883_g N_VDD_Mp8@1883_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1882 N_OUT8_Mp8@1882_d N_OUT7_Mp8@1882_g N_VDD_Mp8@1882_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1881 N_OUT8_Mn8@1881_d N_OUT7_Mn8@1881_g N_VSS_Mn8@1881_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1880 N_OUT8_Mn8@1880_d N_OUT7_Mn8@1880_g N_VSS_Mn8@1880_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1881 N_OUT8_Mp8@1881_d N_OUT7_Mp8@1881_g N_VDD_Mp8@1881_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1880 N_OUT8_Mp8@1880_d N_OUT7_Mp8@1880_g N_VDD_Mp8@1880_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1879 N_OUT8_Mn8@1879_d N_OUT7_Mn8@1879_g N_VSS_Mn8@1879_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1878 N_OUT8_Mn8@1878_d N_OUT7_Mn8@1878_g N_VSS_Mn8@1878_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1879 N_OUT8_Mp8@1879_d N_OUT7_Mp8@1879_g N_VDD_Mp8@1879_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1878 N_OUT8_Mp8@1878_d N_OUT7_Mp8@1878_g N_VDD_Mp8@1878_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1877 N_OUT8_Mn8@1877_d N_OUT7_Mn8@1877_g N_VSS_Mn8@1877_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1876 N_OUT8_Mn8@1876_d N_OUT7_Mn8@1876_g N_VSS_Mn8@1876_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1877 N_OUT8_Mp8@1877_d N_OUT7_Mp8@1877_g N_VDD_Mp8@1877_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1876 N_OUT8_Mp8@1876_d N_OUT7_Mp8@1876_g N_VDD_Mp8@1876_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1875 N_OUT8_Mn8@1875_d N_OUT7_Mn8@1875_g N_VSS_Mn8@1875_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1874 N_OUT8_Mn8@1874_d N_OUT7_Mn8@1874_g N_VSS_Mn8@1874_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1875 N_OUT8_Mp8@1875_d N_OUT7_Mp8@1875_g N_VDD_Mp8@1875_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1874 N_OUT8_Mp8@1874_d N_OUT7_Mp8@1874_g N_VDD_Mp8@1874_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1873 N_OUT8_Mn8@1873_d N_OUT7_Mn8@1873_g N_VSS_Mn8@1873_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1872 N_OUT8_Mn8@1872_d N_OUT7_Mn8@1872_g N_VSS_Mn8@1872_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1873 N_OUT8_Mp8@1873_d N_OUT7_Mp8@1873_g N_VDD_Mp8@1873_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1872 N_OUT8_Mp8@1872_d N_OUT7_Mp8@1872_g N_VDD_Mp8@1872_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1871 N_OUT8_Mn8@1871_d N_OUT7_Mn8@1871_g N_VSS_Mn8@1871_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1870 N_OUT8_Mn8@1870_d N_OUT7_Mn8@1870_g N_VSS_Mn8@1870_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1871 N_OUT8_Mp8@1871_d N_OUT7_Mp8@1871_g N_VDD_Mp8@1871_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1870 N_OUT8_Mp8@1870_d N_OUT7_Mp8@1870_g N_VDD_Mp8@1870_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1869 N_OUT8_Mn8@1869_d N_OUT7_Mn8@1869_g N_VSS_Mn8@1869_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1868 N_OUT8_Mn8@1868_d N_OUT7_Mn8@1868_g N_VSS_Mn8@1868_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1869 N_OUT8_Mp8@1869_d N_OUT7_Mp8@1869_g N_VDD_Mp8@1869_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1868 N_OUT8_Mp8@1868_d N_OUT7_Mp8@1868_g N_VDD_Mp8@1868_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1867 N_OUT8_Mn8@1867_d N_OUT7_Mn8@1867_g N_VSS_Mn8@1867_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1866 N_OUT8_Mn8@1866_d N_OUT7_Mn8@1866_g N_VSS_Mn8@1866_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1867 N_OUT8_Mp8@1867_d N_OUT7_Mp8@1867_g N_VDD_Mp8@1867_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1866 N_OUT8_Mp8@1866_d N_OUT7_Mp8@1866_g N_VDD_Mp8@1866_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1865 N_OUT8_Mn8@1865_d N_OUT7_Mn8@1865_g N_VSS_Mn8@1865_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1864 N_OUT8_Mn8@1864_d N_OUT7_Mn8@1864_g N_VSS_Mn8@1864_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1865 N_OUT8_Mp8@1865_d N_OUT7_Mp8@1865_g N_VDD_Mp8@1865_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1864 N_OUT8_Mp8@1864_d N_OUT7_Mp8@1864_g N_VDD_Mp8@1864_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1863 N_OUT8_Mn8@1863_d N_OUT7_Mn8@1863_g N_VSS_Mn8@1863_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1862 N_OUT8_Mn8@1862_d N_OUT7_Mn8@1862_g N_VSS_Mn8@1862_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1863 N_OUT8_Mp8@1863_d N_OUT7_Mp8@1863_g N_VDD_Mp8@1863_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1862 N_OUT8_Mp8@1862_d N_OUT7_Mp8@1862_g N_VDD_Mp8@1862_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1861 N_OUT8_Mn8@1861_d N_OUT7_Mn8@1861_g N_VSS_Mn8@1861_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1860 N_OUT8_Mn8@1860_d N_OUT7_Mn8@1860_g N_VSS_Mn8@1860_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1861 N_OUT8_Mp8@1861_d N_OUT7_Mp8@1861_g N_VDD_Mp8@1861_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1860 N_OUT8_Mp8@1860_d N_OUT7_Mp8@1860_g N_VDD_Mp8@1860_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1859 N_OUT8_Mn8@1859_d N_OUT7_Mn8@1859_g N_VSS_Mn8@1859_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1858 N_OUT8_Mn8@1858_d N_OUT7_Mn8@1858_g N_VSS_Mn8@1858_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1859 N_OUT8_Mp8@1859_d N_OUT7_Mp8@1859_g N_VDD_Mp8@1859_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1858 N_OUT8_Mp8@1858_d N_OUT7_Mp8@1858_g N_VDD_Mp8@1858_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1857 N_OUT8_Mn8@1857_d N_OUT7_Mn8@1857_g N_VSS_Mn8@1857_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1856 N_OUT8_Mn8@1856_d N_OUT7_Mn8@1856_g N_VSS_Mn8@1856_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1857 N_OUT8_Mp8@1857_d N_OUT7_Mp8@1857_g N_VDD_Mp8@1857_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1856 N_OUT8_Mp8@1856_d N_OUT7_Mp8@1856_g N_VDD_Mp8@1856_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1855 N_OUT8_Mn8@1855_d N_OUT7_Mn8@1855_g N_VSS_Mn8@1855_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1854 N_OUT8_Mn8@1854_d N_OUT7_Mn8@1854_g N_VSS_Mn8@1854_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1855 N_OUT8_Mp8@1855_d N_OUT7_Mp8@1855_g N_VDD_Mp8@1855_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1854 N_OUT8_Mp8@1854_d N_OUT7_Mp8@1854_g N_VDD_Mp8@1854_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1853 N_OUT8_Mn8@1853_d N_OUT7_Mn8@1853_g N_VSS_Mn8@1853_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1852 N_OUT8_Mn8@1852_d N_OUT7_Mn8@1852_g N_VSS_Mn8@1852_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1853 N_OUT8_Mp8@1853_d N_OUT7_Mp8@1853_g N_VDD_Mp8@1853_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1852 N_OUT8_Mp8@1852_d N_OUT7_Mp8@1852_g N_VDD_Mp8@1852_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1851 N_OUT8_Mn8@1851_d N_OUT7_Mn8@1851_g N_VSS_Mn8@1851_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1850 N_OUT8_Mn8@1850_d N_OUT7_Mn8@1850_g N_VSS_Mn8@1850_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1851 N_OUT8_Mp8@1851_d N_OUT7_Mp8@1851_g N_VDD_Mp8@1851_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1850 N_OUT8_Mp8@1850_d N_OUT7_Mp8@1850_g N_VDD_Mp8@1850_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1849 N_OUT8_Mn8@1849_d N_OUT7_Mn8@1849_g N_VSS_Mn8@1849_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1848 N_OUT8_Mn8@1848_d N_OUT7_Mn8@1848_g N_VSS_Mn8@1848_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1849 N_OUT8_Mp8@1849_d N_OUT7_Mp8@1849_g N_VDD_Mp8@1849_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1848 N_OUT8_Mp8@1848_d N_OUT7_Mp8@1848_g N_VDD_Mp8@1848_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1847 N_OUT8_Mn8@1847_d N_OUT7_Mn8@1847_g N_VSS_Mn8@1847_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1846 N_OUT8_Mn8@1846_d N_OUT7_Mn8@1846_g N_VSS_Mn8@1846_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1847 N_OUT8_Mp8@1847_d N_OUT7_Mp8@1847_g N_VDD_Mp8@1847_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1846 N_OUT8_Mp8@1846_d N_OUT7_Mp8@1846_g N_VDD_Mp8@1846_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1845 N_OUT8_Mn8@1845_d N_OUT7_Mn8@1845_g N_VSS_Mn8@1845_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1844 N_OUT8_Mn8@1844_d N_OUT7_Mn8@1844_g N_VSS_Mn8@1844_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1845 N_OUT8_Mp8@1845_d N_OUT7_Mp8@1845_g N_VDD_Mp8@1845_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1844 N_OUT8_Mp8@1844_d N_OUT7_Mp8@1844_g N_VDD_Mp8@1844_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1843 N_OUT8_Mn8@1843_d N_OUT7_Mn8@1843_g N_VSS_Mn8@1843_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1842 N_OUT8_Mn8@1842_d N_OUT7_Mn8@1842_g N_VSS_Mn8@1842_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1843 N_OUT8_Mp8@1843_d N_OUT7_Mp8@1843_g N_VDD_Mp8@1843_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1842 N_OUT8_Mp8@1842_d N_OUT7_Mp8@1842_g N_VDD_Mp8@1842_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1841 N_OUT8_Mn8@1841_d N_OUT7_Mn8@1841_g N_VSS_Mn8@1841_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1840 N_OUT8_Mn8@1840_d N_OUT7_Mn8@1840_g N_VSS_Mn8@1840_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1841 N_OUT8_Mp8@1841_d N_OUT7_Mp8@1841_g N_VDD_Mp8@1841_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1840 N_OUT8_Mp8@1840_d N_OUT7_Mp8@1840_g N_VDD_Mp8@1840_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1839 N_OUT8_Mn8@1839_d N_OUT7_Mn8@1839_g N_VSS_Mn8@1839_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1838 N_OUT8_Mn8@1838_d N_OUT7_Mn8@1838_g N_VSS_Mn8@1838_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1839 N_OUT8_Mp8@1839_d N_OUT7_Mp8@1839_g N_VDD_Mp8@1839_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1838 N_OUT8_Mp8@1838_d N_OUT7_Mp8@1838_g N_VDD_Mp8@1838_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1837 N_OUT8_Mn8@1837_d N_OUT7_Mn8@1837_g N_VSS_Mn8@1837_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1836 N_OUT8_Mn8@1836_d N_OUT7_Mn8@1836_g N_VSS_Mn8@1836_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1837 N_OUT8_Mp8@1837_d N_OUT7_Mp8@1837_g N_VDD_Mp8@1837_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1836 N_OUT8_Mp8@1836_d N_OUT7_Mp8@1836_g N_VDD_Mp8@1836_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1835 N_OUT8_Mn8@1835_d N_OUT7_Mn8@1835_g N_VSS_Mn8@1835_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1834 N_OUT8_Mn8@1834_d N_OUT7_Mn8@1834_g N_VSS_Mn8@1834_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1835 N_OUT8_Mp8@1835_d N_OUT7_Mp8@1835_g N_VDD_Mp8@1835_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1834 N_OUT8_Mp8@1834_d N_OUT7_Mp8@1834_g N_VDD_Mp8@1834_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1833 N_OUT8_Mn8@1833_d N_OUT7_Mn8@1833_g N_VSS_Mn8@1833_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1832 N_OUT8_Mn8@1832_d N_OUT7_Mn8@1832_g N_VSS_Mn8@1832_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1833 N_OUT8_Mp8@1833_d N_OUT7_Mp8@1833_g N_VDD_Mp8@1833_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1832 N_OUT8_Mp8@1832_d N_OUT7_Mp8@1832_g N_VDD_Mp8@1832_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1831 N_OUT8_Mn8@1831_d N_OUT7_Mn8@1831_g N_VSS_Mn8@1831_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1830 N_OUT8_Mn8@1830_d N_OUT7_Mn8@1830_g N_VSS_Mn8@1830_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1831 N_OUT8_Mp8@1831_d N_OUT7_Mp8@1831_g N_VDD_Mp8@1831_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1830 N_OUT8_Mp8@1830_d N_OUT7_Mp8@1830_g N_VDD_Mp8@1830_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1829 N_OUT8_Mn8@1829_d N_OUT7_Mn8@1829_g N_VSS_Mn8@1829_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1828 N_OUT8_Mn8@1828_d N_OUT7_Mn8@1828_g N_VSS_Mn8@1828_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1829 N_OUT8_Mp8@1829_d N_OUT7_Mp8@1829_g N_VDD_Mp8@1829_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1828 N_OUT8_Mp8@1828_d N_OUT7_Mp8@1828_g N_VDD_Mp8@1828_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1827 N_OUT8_Mn8@1827_d N_OUT7_Mn8@1827_g N_VSS_Mn8@1827_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1826 N_OUT8_Mn8@1826_d N_OUT7_Mn8@1826_g N_VSS_Mn8@1826_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1827 N_OUT8_Mp8@1827_d N_OUT7_Mp8@1827_g N_VDD_Mp8@1827_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1826 N_OUT8_Mp8@1826_d N_OUT7_Mp8@1826_g N_VDD_Mp8@1826_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1825 N_OUT8_Mn8@1825_d N_OUT7_Mn8@1825_g N_VSS_Mn8@1825_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1824 N_OUT8_Mn8@1824_d N_OUT7_Mn8@1824_g N_VSS_Mn8@1824_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1825 N_OUT8_Mp8@1825_d N_OUT7_Mp8@1825_g N_VDD_Mp8@1825_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1824 N_OUT8_Mp8@1824_d N_OUT7_Mp8@1824_g N_VDD_Mp8@1824_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1823 N_OUT8_Mn8@1823_d N_OUT7_Mn8@1823_g N_VSS_Mn8@1823_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1822 N_OUT8_Mn8@1822_d N_OUT7_Mn8@1822_g N_VSS_Mn8@1822_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1823 N_OUT8_Mp8@1823_d N_OUT7_Mp8@1823_g N_VDD_Mp8@1823_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1822 N_OUT8_Mp8@1822_d N_OUT7_Mp8@1822_g N_VDD_Mp8@1822_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1821 N_OUT8_Mn8@1821_d N_OUT7_Mn8@1821_g N_VSS_Mn8@1821_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1820 N_OUT8_Mn8@1820_d N_OUT7_Mn8@1820_g N_VSS_Mn8@1820_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1821 N_OUT8_Mp8@1821_d N_OUT7_Mp8@1821_g N_VDD_Mp8@1821_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1820 N_OUT8_Mp8@1820_d N_OUT7_Mp8@1820_g N_VDD_Mp8@1820_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1819 N_OUT8_Mn8@1819_d N_OUT7_Mn8@1819_g N_VSS_Mn8@1819_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1818 N_OUT8_Mn8@1818_d N_OUT7_Mn8@1818_g N_VSS_Mn8@1818_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1819 N_OUT8_Mp8@1819_d N_OUT7_Mp8@1819_g N_VDD_Mp8@1819_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1818 N_OUT8_Mp8@1818_d N_OUT7_Mp8@1818_g N_VDD_Mp8@1818_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1817 N_OUT8_Mn8@1817_d N_OUT7_Mn8@1817_g N_VSS_Mn8@1817_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1816 N_OUT8_Mn8@1816_d N_OUT7_Mn8@1816_g N_VSS_Mn8@1816_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1817 N_OUT8_Mp8@1817_d N_OUT7_Mp8@1817_g N_VDD_Mp8@1817_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1816 N_OUT8_Mp8@1816_d N_OUT7_Mp8@1816_g N_VDD_Mp8@1816_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1815 N_OUT8_Mn8@1815_d N_OUT7_Mn8@1815_g N_VSS_Mn8@1815_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1814 N_OUT8_Mn8@1814_d N_OUT7_Mn8@1814_g N_VSS_Mn8@1814_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1815 N_OUT8_Mp8@1815_d N_OUT7_Mp8@1815_g N_VDD_Mp8@1815_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1814 N_OUT8_Mp8@1814_d N_OUT7_Mp8@1814_g N_VDD_Mp8@1814_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1813 N_OUT8_Mn8@1813_d N_OUT7_Mn8@1813_g N_VSS_Mn8@1813_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1812 N_OUT8_Mn8@1812_d N_OUT7_Mn8@1812_g N_VSS_Mn8@1812_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1813 N_OUT8_Mp8@1813_d N_OUT7_Mp8@1813_g N_VDD_Mp8@1813_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1812 N_OUT8_Mp8@1812_d N_OUT7_Mp8@1812_g N_VDD_Mp8@1812_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1811 N_OUT8_Mn8@1811_d N_OUT7_Mn8@1811_g N_VSS_Mn8@1811_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1810 N_OUT8_Mn8@1810_d N_OUT7_Mn8@1810_g N_VSS_Mn8@1810_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1811 N_OUT8_Mp8@1811_d N_OUT7_Mp8@1811_g N_VDD_Mp8@1811_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1810 N_OUT8_Mp8@1810_d N_OUT7_Mp8@1810_g N_VDD_Mp8@1810_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1809 N_OUT8_Mn8@1809_d N_OUT7_Mn8@1809_g N_VSS_Mn8@1809_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1808 N_OUT8_Mn8@1808_d N_OUT7_Mn8@1808_g N_VSS_Mn8@1808_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1809 N_OUT8_Mp8@1809_d N_OUT7_Mp8@1809_g N_VDD_Mp8@1809_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1808 N_OUT8_Mp8@1808_d N_OUT7_Mp8@1808_g N_VDD_Mp8@1808_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1807 N_OUT8_Mn8@1807_d N_OUT7_Mn8@1807_g N_VSS_Mn8@1807_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1806 N_OUT8_Mn8@1806_d N_OUT7_Mn8@1806_g N_VSS_Mn8@1806_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1807 N_OUT8_Mp8@1807_d N_OUT7_Mp8@1807_g N_VDD_Mp8@1807_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1806 N_OUT8_Mp8@1806_d N_OUT7_Mp8@1806_g N_VDD_Mp8@1806_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1805 N_OUT8_Mn8@1805_d N_OUT7_Mn8@1805_g N_VSS_Mn8@1805_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1804 N_OUT8_Mn8@1804_d N_OUT7_Mn8@1804_g N_VSS_Mn8@1804_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1805 N_OUT8_Mp8@1805_d N_OUT7_Mp8@1805_g N_VDD_Mp8@1805_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1804 N_OUT8_Mp8@1804_d N_OUT7_Mp8@1804_g N_VDD_Mp8@1804_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1803 N_OUT8_Mn8@1803_d N_OUT7_Mn8@1803_g N_VSS_Mn8@1803_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1802 N_OUT8_Mn8@1802_d N_OUT7_Mn8@1802_g N_VSS_Mn8@1802_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1803 N_OUT8_Mp8@1803_d N_OUT7_Mp8@1803_g N_VDD_Mp8@1803_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1802 N_OUT8_Mp8@1802_d N_OUT7_Mp8@1802_g N_VDD_Mp8@1802_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1801 N_OUT8_Mn8@1801_d N_OUT7_Mn8@1801_g N_VSS_Mn8@1801_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1800 N_OUT8_Mn8@1800_d N_OUT7_Mn8@1800_g N_VSS_Mn8@1800_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1801 N_OUT8_Mp8@1801_d N_OUT7_Mp8@1801_g N_VDD_Mp8@1801_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1800 N_OUT8_Mp8@1800_d N_OUT7_Mp8@1800_g N_VDD_Mp8@1800_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1799 N_OUT8_Mn8@1799_d N_OUT7_Mn8@1799_g N_VSS_Mn8@1799_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1798 N_OUT8_Mn8@1798_d N_OUT7_Mn8@1798_g N_VSS_Mn8@1798_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1799 N_OUT8_Mp8@1799_d N_OUT7_Mp8@1799_g N_VDD_Mp8@1799_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1798 N_OUT8_Mp8@1798_d N_OUT7_Mp8@1798_g N_VDD_Mp8@1798_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1797 N_OUT8_Mn8@1797_d N_OUT7_Mn8@1797_g N_VSS_Mn8@1797_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1796 N_OUT8_Mn8@1796_d N_OUT7_Mn8@1796_g N_VSS_Mn8@1796_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1797 N_OUT8_Mp8@1797_d N_OUT7_Mp8@1797_g N_VDD_Mp8@1797_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1796 N_OUT8_Mp8@1796_d N_OUT7_Mp8@1796_g N_VDD_Mp8@1796_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1795 N_OUT8_Mn8@1795_d N_OUT7_Mn8@1795_g N_VSS_Mn8@1795_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1794 N_OUT8_Mn8@1794_d N_OUT7_Mn8@1794_g N_VSS_Mn8@1794_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1795 N_OUT8_Mp8@1795_d N_OUT7_Mp8@1795_g N_VDD_Mp8@1795_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1794 N_OUT8_Mp8@1794_d N_OUT7_Mp8@1794_g N_VDD_Mp8@1794_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1793 N_OUT8_Mn8@1793_d N_OUT7_Mn8@1793_g N_VSS_Mn8@1793_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1792 N_OUT8_Mn8@1792_d N_OUT7_Mn8@1792_g N_VSS_Mn8@1792_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1793 N_OUT8_Mp8@1793_d N_OUT7_Mp8@1793_g N_VDD_Mp8@1793_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1792 N_OUT8_Mp8@1792_d N_OUT7_Mp8@1792_g N_VDD_Mp8@1792_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1791 N_OUT8_Mn8@1791_d N_OUT7_Mn8@1791_g N_VSS_Mn8@1791_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1790 N_OUT8_Mn8@1790_d N_OUT7_Mn8@1790_g N_VSS_Mn8@1790_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1791 N_OUT8_Mp8@1791_d N_OUT7_Mp8@1791_g N_VDD_Mp8@1791_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1790 N_OUT8_Mp8@1790_d N_OUT7_Mp8@1790_g N_VDD_Mp8@1790_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1789 N_OUT8_Mn8@1789_d N_OUT7_Mn8@1789_g N_VSS_Mn8@1789_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1788 N_OUT8_Mn8@1788_d N_OUT7_Mn8@1788_g N_VSS_Mn8@1788_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1789 N_OUT8_Mp8@1789_d N_OUT7_Mp8@1789_g N_VDD_Mp8@1789_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1788 N_OUT8_Mp8@1788_d N_OUT7_Mp8@1788_g N_VDD_Mp8@1788_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1787 N_OUT8_Mn8@1787_d N_OUT7_Mn8@1787_g N_VSS_Mn8@1787_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1786 N_OUT8_Mn8@1786_d N_OUT7_Mn8@1786_g N_VSS_Mn8@1786_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1787 N_OUT8_Mp8@1787_d N_OUT7_Mp8@1787_g N_VDD_Mp8@1787_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1786 N_OUT8_Mp8@1786_d N_OUT7_Mp8@1786_g N_VDD_Mp8@1786_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1785 N_OUT8_Mn8@1785_d N_OUT7_Mn8@1785_g N_VSS_Mn8@1785_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1784 N_OUT8_Mn8@1784_d N_OUT7_Mn8@1784_g N_VSS_Mn8@1784_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1785 N_OUT8_Mp8@1785_d N_OUT7_Mp8@1785_g N_VDD_Mp8@1785_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1784 N_OUT8_Mp8@1784_d N_OUT7_Mp8@1784_g N_VDD_Mp8@1784_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1783 N_OUT8_Mn8@1783_d N_OUT7_Mn8@1783_g N_VSS_Mn8@1783_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1782 N_OUT8_Mn8@1782_d N_OUT7_Mn8@1782_g N_VSS_Mn8@1782_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1783 N_OUT8_Mp8@1783_d N_OUT7_Mp8@1783_g N_VDD_Mp8@1783_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1782 N_OUT8_Mp8@1782_d N_OUT7_Mp8@1782_g N_VDD_Mp8@1782_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1781 N_OUT8_Mn8@1781_d N_OUT7_Mn8@1781_g N_VSS_Mn8@1781_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1780 N_OUT8_Mn8@1780_d N_OUT7_Mn8@1780_g N_VSS_Mn8@1780_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1781 N_OUT8_Mp8@1781_d N_OUT7_Mp8@1781_g N_VDD_Mp8@1781_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1780 N_OUT8_Mp8@1780_d N_OUT7_Mp8@1780_g N_VDD_Mp8@1780_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1779 N_OUT8_Mn8@1779_d N_OUT7_Mn8@1779_g N_VSS_Mn8@1779_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1778 N_OUT8_Mn8@1778_d N_OUT7_Mn8@1778_g N_VSS_Mn8@1778_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1779 N_OUT8_Mp8@1779_d N_OUT7_Mp8@1779_g N_VDD_Mp8@1779_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1778 N_OUT8_Mp8@1778_d N_OUT7_Mp8@1778_g N_VDD_Mp8@1778_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1777 N_OUT8_Mn8@1777_d N_OUT7_Mn8@1777_g N_VSS_Mn8@1777_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1776 N_OUT8_Mn8@1776_d N_OUT7_Mn8@1776_g N_VSS_Mn8@1776_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1777 N_OUT8_Mp8@1777_d N_OUT7_Mp8@1777_g N_VDD_Mp8@1777_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1776 N_OUT8_Mp8@1776_d N_OUT7_Mp8@1776_g N_VDD_Mp8@1776_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1775 N_OUT8_Mn8@1775_d N_OUT7_Mn8@1775_g N_VSS_Mn8@1775_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1774 N_OUT8_Mn8@1774_d N_OUT7_Mn8@1774_g N_VSS_Mn8@1774_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1775 N_OUT8_Mp8@1775_d N_OUT7_Mp8@1775_g N_VDD_Mp8@1775_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1774 N_OUT8_Mp8@1774_d N_OUT7_Mp8@1774_g N_VDD_Mp8@1774_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1773 N_OUT8_Mn8@1773_d N_OUT7_Mn8@1773_g N_VSS_Mn8@1773_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1772 N_OUT8_Mn8@1772_d N_OUT7_Mn8@1772_g N_VSS_Mn8@1772_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1773 N_OUT8_Mp8@1773_d N_OUT7_Mp8@1773_g N_VDD_Mp8@1773_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1772 N_OUT8_Mp8@1772_d N_OUT7_Mp8@1772_g N_VDD_Mp8@1772_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1771 N_OUT8_Mn8@1771_d N_OUT7_Mn8@1771_g N_VSS_Mn8@1771_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1770 N_OUT8_Mn8@1770_d N_OUT7_Mn8@1770_g N_VSS_Mn8@1770_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1771 N_OUT8_Mp8@1771_d N_OUT7_Mp8@1771_g N_VDD_Mp8@1771_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1770 N_OUT8_Mp8@1770_d N_OUT7_Mp8@1770_g N_VDD_Mp8@1770_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1769 N_OUT8_Mn8@1769_d N_OUT7_Mn8@1769_g N_VSS_Mn8@1769_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1768 N_OUT8_Mn8@1768_d N_OUT7_Mn8@1768_g N_VSS_Mn8@1768_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1769 N_OUT8_Mp8@1769_d N_OUT7_Mp8@1769_g N_VDD_Mp8@1769_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1768 N_OUT8_Mp8@1768_d N_OUT7_Mp8@1768_g N_VDD_Mp8@1768_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1767 N_OUT8_Mn8@1767_d N_OUT7_Mn8@1767_g N_VSS_Mn8@1767_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1766 N_OUT8_Mn8@1766_d N_OUT7_Mn8@1766_g N_VSS_Mn8@1766_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1767 N_OUT8_Mp8@1767_d N_OUT7_Mp8@1767_g N_VDD_Mp8@1767_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1766 N_OUT8_Mp8@1766_d N_OUT7_Mp8@1766_g N_VDD_Mp8@1766_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1765 N_OUT8_Mn8@1765_d N_OUT7_Mn8@1765_g N_VSS_Mn8@1765_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1764 N_OUT8_Mn8@1764_d N_OUT7_Mn8@1764_g N_VSS_Mn8@1764_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1765 N_OUT8_Mp8@1765_d N_OUT7_Mp8@1765_g N_VDD_Mp8@1765_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1764 N_OUT8_Mp8@1764_d N_OUT7_Mp8@1764_g N_VDD_Mp8@1764_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1763 N_OUT8_Mn8@1763_d N_OUT7_Mn8@1763_g N_VSS_Mn8@1763_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1762 N_OUT8_Mn8@1762_d N_OUT7_Mn8@1762_g N_VSS_Mn8@1762_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1763 N_OUT8_Mp8@1763_d N_OUT7_Mp8@1763_g N_VDD_Mp8@1763_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1762 N_OUT8_Mp8@1762_d N_OUT7_Mp8@1762_g N_VDD_Mp8@1762_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1761 N_OUT8_Mn8@1761_d N_OUT7_Mn8@1761_g N_VSS_Mn8@1761_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1760 N_OUT8_Mn8@1760_d N_OUT7_Mn8@1760_g N_VSS_Mn8@1760_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1761 N_OUT8_Mp8@1761_d N_OUT7_Mp8@1761_g N_VDD_Mp8@1761_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1760 N_OUT8_Mp8@1760_d N_OUT7_Mp8@1760_g N_VDD_Mp8@1760_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1759 N_OUT8_Mn8@1759_d N_OUT7_Mn8@1759_g N_VSS_Mn8@1759_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1758 N_OUT8_Mn8@1758_d N_OUT7_Mn8@1758_g N_VSS_Mn8@1758_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1759 N_OUT8_Mp8@1759_d N_OUT7_Mp8@1759_g N_VDD_Mp8@1759_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1758 N_OUT8_Mp8@1758_d N_OUT7_Mp8@1758_g N_VDD_Mp8@1758_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1757 N_OUT8_Mn8@1757_d N_OUT7_Mn8@1757_g N_VSS_Mn8@1757_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1756 N_OUT8_Mn8@1756_d N_OUT7_Mn8@1756_g N_VSS_Mn8@1756_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1757 N_OUT8_Mp8@1757_d N_OUT7_Mp8@1757_g N_VDD_Mp8@1757_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1756 N_OUT8_Mp8@1756_d N_OUT7_Mp8@1756_g N_VDD_Mp8@1756_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1755 N_OUT8_Mn8@1755_d N_OUT7_Mn8@1755_g N_VSS_Mn8@1755_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1754 N_OUT8_Mn8@1754_d N_OUT7_Mn8@1754_g N_VSS_Mn8@1754_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1755 N_OUT8_Mp8@1755_d N_OUT7_Mp8@1755_g N_VDD_Mp8@1755_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1754 N_OUT8_Mp8@1754_d N_OUT7_Mp8@1754_g N_VDD_Mp8@1754_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1753 N_OUT8_Mn8@1753_d N_OUT7_Mn8@1753_g N_VSS_Mn8@1753_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1752 N_OUT8_Mn8@1752_d N_OUT7_Mn8@1752_g N_VSS_Mn8@1752_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1753 N_OUT8_Mp8@1753_d N_OUT7_Mp8@1753_g N_VDD_Mp8@1753_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1752 N_OUT8_Mp8@1752_d N_OUT7_Mp8@1752_g N_VDD_Mp8@1752_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1751 N_OUT8_Mn8@1751_d N_OUT7_Mn8@1751_g N_VSS_Mn8@1751_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1750 N_OUT8_Mn8@1750_d N_OUT7_Mn8@1750_g N_VSS_Mn8@1750_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1751 N_OUT8_Mp8@1751_d N_OUT7_Mp8@1751_g N_VDD_Mp8@1751_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1750 N_OUT8_Mp8@1750_d N_OUT7_Mp8@1750_g N_VDD_Mp8@1750_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1749 N_OUT8_Mn8@1749_d N_OUT7_Mn8@1749_g N_VSS_Mn8@1749_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1748 N_OUT8_Mn8@1748_d N_OUT7_Mn8@1748_g N_VSS_Mn8@1748_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1749 N_OUT8_Mp8@1749_d N_OUT7_Mp8@1749_g N_VDD_Mp8@1749_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1748 N_OUT8_Mp8@1748_d N_OUT7_Mp8@1748_g N_VDD_Mp8@1748_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1747 N_OUT8_Mn8@1747_d N_OUT7_Mn8@1747_g N_VSS_Mn8@1747_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1746 N_OUT8_Mn8@1746_d N_OUT7_Mn8@1746_g N_VSS_Mn8@1746_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1747 N_OUT8_Mp8@1747_d N_OUT7_Mp8@1747_g N_VDD_Mp8@1747_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1746 N_OUT8_Mp8@1746_d N_OUT7_Mp8@1746_g N_VDD_Mp8@1746_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1745 N_OUT8_Mn8@1745_d N_OUT7_Mn8@1745_g N_VSS_Mn8@1745_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1744 N_OUT8_Mn8@1744_d N_OUT7_Mn8@1744_g N_VSS_Mn8@1744_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1745 N_OUT8_Mp8@1745_d N_OUT7_Mp8@1745_g N_VDD_Mp8@1745_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1744 N_OUT8_Mp8@1744_d N_OUT7_Mp8@1744_g N_VDD_Mp8@1744_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1743 N_OUT8_Mn8@1743_d N_OUT7_Mn8@1743_g N_VSS_Mn8@1743_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1742 N_OUT8_Mn8@1742_d N_OUT7_Mn8@1742_g N_VSS_Mn8@1742_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1743 N_OUT8_Mp8@1743_d N_OUT7_Mp8@1743_g N_VDD_Mp8@1743_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1742 N_OUT8_Mp8@1742_d N_OUT7_Mp8@1742_g N_VDD_Mp8@1742_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1741 N_OUT8_Mn8@1741_d N_OUT7_Mn8@1741_g N_VSS_Mn8@1741_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1740 N_OUT8_Mn8@1740_d N_OUT7_Mn8@1740_g N_VSS_Mn8@1740_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1741 N_OUT8_Mp8@1741_d N_OUT7_Mp8@1741_g N_VDD_Mp8@1741_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1740 N_OUT8_Mp8@1740_d N_OUT7_Mp8@1740_g N_VDD_Mp8@1740_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1739 N_OUT8_Mn8@1739_d N_OUT7_Mn8@1739_g N_VSS_Mn8@1739_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1738 N_OUT8_Mn8@1738_d N_OUT7_Mn8@1738_g N_VSS_Mn8@1738_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1739 N_OUT8_Mp8@1739_d N_OUT7_Mp8@1739_g N_VDD_Mp8@1739_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1738 N_OUT8_Mp8@1738_d N_OUT7_Mp8@1738_g N_VDD_Mp8@1738_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1737 N_OUT8_Mn8@1737_d N_OUT7_Mn8@1737_g N_VSS_Mn8@1737_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1736 N_OUT8_Mn8@1736_d N_OUT7_Mn8@1736_g N_VSS_Mn8@1736_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1737 N_OUT8_Mp8@1737_d N_OUT7_Mp8@1737_g N_VDD_Mp8@1737_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1736 N_OUT8_Mp8@1736_d N_OUT7_Mp8@1736_g N_VDD_Mp8@1736_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1735 N_OUT8_Mn8@1735_d N_OUT7_Mn8@1735_g N_VSS_Mn8@1735_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1734 N_OUT8_Mn8@1734_d N_OUT7_Mn8@1734_g N_VSS_Mn8@1734_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1735 N_OUT8_Mp8@1735_d N_OUT7_Mp8@1735_g N_VDD_Mp8@1735_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1734 N_OUT8_Mp8@1734_d N_OUT7_Mp8@1734_g N_VDD_Mp8@1734_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1733 N_OUT8_Mn8@1733_d N_OUT7_Mn8@1733_g N_VSS_Mn8@1733_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1732 N_OUT8_Mn8@1732_d N_OUT7_Mn8@1732_g N_VSS_Mn8@1732_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1733 N_OUT8_Mp8@1733_d N_OUT7_Mp8@1733_g N_VDD_Mp8@1733_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1732 N_OUT8_Mp8@1732_d N_OUT7_Mp8@1732_g N_VDD_Mp8@1732_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1731 N_OUT8_Mn8@1731_d N_OUT7_Mn8@1731_g N_VSS_Mn8@1731_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1730 N_OUT8_Mn8@1730_d N_OUT7_Mn8@1730_g N_VSS_Mn8@1730_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1731 N_OUT8_Mp8@1731_d N_OUT7_Mp8@1731_g N_VDD_Mp8@1731_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1730 N_OUT8_Mp8@1730_d N_OUT7_Mp8@1730_g N_VDD_Mp8@1730_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1729 N_OUT8_Mn8@1729_d N_OUT7_Mn8@1729_g N_VSS_Mn8@1729_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1728 N_OUT8_Mn8@1728_d N_OUT7_Mn8@1728_g N_VSS_Mn8@1728_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1729 N_OUT8_Mp8@1729_d N_OUT7_Mp8@1729_g N_VDD_Mp8@1729_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1728 N_OUT8_Mp8@1728_d N_OUT7_Mp8@1728_g N_VDD_Mp8@1728_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1727 N_OUT8_Mn8@1727_d N_OUT7_Mn8@1727_g N_VSS_Mn8@1727_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1726 N_OUT8_Mn8@1726_d N_OUT7_Mn8@1726_g N_VSS_Mn8@1726_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1727 N_OUT8_Mp8@1727_d N_OUT7_Mp8@1727_g N_VDD_Mp8@1727_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1726 N_OUT8_Mp8@1726_d N_OUT7_Mp8@1726_g N_VDD_Mp8@1726_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1725 N_OUT8_Mn8@1725_d N_OUT7_Mn8@1725_g N_VSS_Mn8@1725_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1724 N_OUT8_Mn8@1724_d N_OUT7_Mn8@1724_g N_VSS_Mn8@1724_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1725 N_OUT8_Mp8@1725_d N_OUT7_Mp8@1725_g N_VDD_Mp8@1725_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1724 N_OUT8_Mp8@1724_d N_OUT7_Mp8@1724_g N_VDD_Mp8@1724_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1723 N_OUT8_Mn8@1723_d N_OUT7_Mn8@1723_g N_VSS_Mn8@1723_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1722 N_OUT8_Mn8@1722_d N_OUT7_Mn8@1722_g N_VSS_Mn8@1722_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1723 N_OUT8_Mp8@1723_d N_OUT7_Mp8@1723_g N_VDD_Mp8@1723_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1722 N_OUT8_Mp8@1722_d N_OUT7_Mp8@1722_g N_VDD_Mp8@1722_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1721 N_OUT8_Mn8@1721_d N_OUT7_Mn8@1721_g N_VSS_Mn8@1721_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1720 N_OUT8_Mn8@1720_d N_OUT7_Mn8@1720_g N_VSS_Mn8@1720_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1721 N_OUT8_Mp8@1721_d N_OUT7_Mp8@1721_g N_VDD_Mp8@1721_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1720 N_OUT8_Mp8@1720_d N_OUT7_Mp8@1720_g N_VDD_Mp8@1720_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1719 N_OUT8_Mn8@1719_d N_OUT7_Mn8@1719_g N_VSS_Mn8@1719_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1718 N_OUT8_Mn8@1718_d N_OUT7_Mn8@1718_g N_VSS_Mn8@1718_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1719 N_OUT8_Mp8@1719_d N_OUT7_Mp8@1719_g N_VDD_Mp8@1719_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1718 N_OUT8_Mp8@1718_d N_OUT7_Mp8@1718_g N_VDD_Mp8@1718_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1717 N_OUT8_Mn8@1717_d N_OUT7_Mn8@1717_g N_VSS_Mn8@1717_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1716 N_OUT8_Mn8@1716_d N_OUT7_Mn8@1716_g N_VSS_Mn8@1716_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1717 N_OUT8_Mp8@1717_d N_OUT7_Mp8@1717_g N_VDD_Mp8@1717_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1716 N_OUT8_Mp8@1716_d N_OUT7_Mp8@1716_g N_VDD_Mp8@1716_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1715 N_OUT8_Mn8@1715_d N_OUT7_Mn8@1715_g N_VSS_Mn8@1715_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1714 N_OUT8_Mn8@1714_d N_OUT7_Mn8@1714_g N_VSS_Mn8@1714_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1715 N_OUT8_Mp8@1715_d N_OUT7_Mp8@1715_g N_VDD_Mp8@1715_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1714 N_OUT8_Mp8@1714_d N_OUT7_Mp8@1714_g N_VDD_Mp8@1714_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1713 N_OUT8_Mn8@1713_d N_OUT7_Mn8@1713_g N_VSS_Mn8@1713_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1712 N_OUT8_Mn8@1712_d N_OUT7_Mn8@1712_g N_VSS_Mn8@1712_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1713 N_OUT8_Mp8@1713_d N_OUT7_Mp8@1713_g N_VDD_Mp8@1713_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1712 N_OUT8_Mp8@1712_d N_OUT7_Mp8@1712_g N_VDD_Mp8@1712_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1711 N_OUT8_Mn8@1711_d N_OUT7_Mn8@1711_g N_VSS_Mn8@1711_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1710 N_OUT8_Mn8@1710_d N_OUT7_Mn8@1710_g N_VSS_Mn8@1710_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1711 N_OUT8_Mp8@1711_d N_OUT7_Mp8@1711_g N_VDD_Mp8@1711_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1710 N_OUT8_Mp8@1710_d N_OUT7_Mp8@1710_g N_VDD_Mp8@1710_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1709 N_OUT8_Mn8@1709_d N_OUT7_Mn8@1709_g N_VSS_Mn8@1709_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1708 N_OUT8_Mn8@1708_d N_OUT7_Mn8@1708_g N_VSS_Mn8@1708_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1709 N_OUT8_Mp8@1709_d N_OUT7_Mp8@1709_g N_VDD_Mp8@1709_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1708 N_OUT8_Mp8@1708_d N_OUT7_Mp8@1708_g N_VDD_Mp8@1708_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1707 N_OUT8_Mn8@1707_d N_OUT7_Mn8@1707_g N_VSS_Mn8@1707_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1706 N_OUT8_Mn8@1706_d N_OUT7_Mn8@1706_g N_VSS_Mn8@1706_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1707 N_OUT8_Mp8@1707_d N_OUT7_Mp8@1707_g N_VDD_Mp8@1707_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1706 N_OUT8_Mp8@1706_d N_OUT7_Mp8@1706_g N_VDD_Mp8@1706_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1705 N_OUT8_Mn8@1705_d N_OUT7_Mn8@1705_g N_VSS_Mn8@1705_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1704 N_OUT8_Mn8@1704_d N_OUT7_Mn8@1704_g N_VSS_Mn8@1704_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1705 N_OUT8_Mp8@1705_d N_OUT7_Mp8@1705_g N_VDD_Mp8@1705_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1704 N_OUT8_Mp8@1704_d N_OUT7_Mp8@1704_g N_VDD_Mp8@1704_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1703 N_OUT8_Mn8@1703_d N_OUT7_Mn8@1703_g N_VSS_Mn8@1703_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1702 N_OUT8_Mn8@1702_d N_OUT7_Mn8@1702_g N_VSS_Mn8@1702_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1703 N_OUT8_Mp8@1703_d N_OUT7_Mp8@1703_g N_VDD_Mp8@1703_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1702 N_OUT8_Mp8@1702_d N_OUT7_Mp8@1702_g N_VDD_Mp8@1702_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1701 N_OUT8_Mn8@1701_d N_OUT7_Mn8@1701_g N_VSS_Mn8@1701_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1700 N_OUT8_Mn8@1700_d N_OUT7_Mn8@1700_g N_VSS_Mn8@1700_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1701 N_OUT8_Mp8@1701_d N_OUT7_Mp8@1701_g N_VDD_Mp8@1701_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1700 N_OUT8_Mp8@1700_d N_OUT7_Mp8@1700_g N_VDD_Mp8@1700_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1699 N_OUT8_Mn8@1699_d N_OUT7_Mn8@1699_g N_VSS_Mn8@1699_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1698 N_OUT8_Mn8@1698_d N_OUT7_Mn8@1698_g N_VSS_Mn8@1698_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1699 N_OUT8_Mp8@1699_d N_OUT7_Mp8@1699_g N_VDD_Mp8@1699_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1698 N_OUT8_Mp8@1698_d N_OUT7_Mp8@1698_g N_VDD_Mp8@1698_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1697 N_OUT8_Mn8@1697_d N_OUT7_Mn8@1697_g N_VSS_Mn8@1697_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1696 N_OUT8_Mn8@1696_d N_OUT7_Mn8@1696_g N_VSS_Mn8@1696_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1697 N_OUT8_Mp8@1697_d N_OUT7_Mp8@1697_g N_VDD_Mp8@1697_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1696 N_OUT8_Mp8@1696_d N_OUT7_Mp8@1696_g N_VDD_Mp8@1696_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1695 N_OUT8_Mn8@1695_d N_OUT7_Mn8@1695_g N_VSS_Mn8@1695_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1694 N_OUT8_Mn8@1694_d N_OUT7_Mn8@1694_g N_VSS_Mn8@1694_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1695 N_OUT8_Mp8@1695_d N_OUT7_Mp8@1695_g N_VDD_Mp8@1695_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1694 N_OUT8_Mp8@1694_d N_OUT7_Mp8@1694_g N_VDD_Mp8@1694_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1693 N_OUT8_Mn8@1693_d N_OUT7_Mn8@1693_g N_VSS_Mn8@1693_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1692 N_OUT8_Mn8@1692_d N_OUT7_Mn8@1692_g N_VSS_Mn8@1692_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1693 N_OUT8_Mp8@1693_d N_OUT7_Mp8@1693_g N_VDD_Mp8@1693_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1692 N_OUT8_Mp8@1692_d N_OUT7_Mp8@1692_g N_VDD_Mp8@1692_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1691 N_OUT8_Mn8@1691_d N_OUT7_Mn8@1691_g N_VSS_Mn8@1691_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1690 N_OUT8_Mn8@1690_d N_OUT7_Mn8@1690_g N_VSS_Mn8@1690_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1691 N_OUT8_Mp8@1691_d N_OUT7_Mp8@1691_g N_VDD_Mp8@1691_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1690 N_OUT8_Mp8@1690_d N_OUT7_Mp8@1690_g N_VDD_Mp8@1690_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1689 N_OUT8_Mn8@1689_d N_OUT7_Mn8@1689_g N_VSS_Mn8@1689_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1688 N_OUT8_Mn8@1688_d N_OUT7_Mn8@1688_g N_VSS_Mn8@1688_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1689 N_OUT8_Mp8@1689_d N_OUT7_Mp8@1689_g N_VDD_Mp8@1689_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1688 N_OUT8_Mp8@1688_d N_OUT7_Mp8@1688_g N_VDD_Mp8@1688_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1687 N_OUT8_Mn8@1687_d N_OUT7_Mn8@1687_g N_VSS_Mn8@1687_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1686 N_OUT8_Mn8@1686_d N_OUT7_Mn8@1686_g N_VSS_Mn8@1686_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1687 N_OUT8_Mp8@1687_d N_OUT7_Mp8@1687_g N_VDD_Mp8@1687_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1686 N_OUT8_Mp8@1686_d N_OUT7_Mp8@1686_g N_VDD_Mp8@1686_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1685 N_OUT8_Mn8@1685_d N_OUT7_Mn8@1685_g N_VSS_Mn8@1685_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1684 N_OUT8_Mn8@1684_d N_OUT7_Mn8@1684_g N_VSS_Mn8@1684_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1685 N_OUT8_Mp8@1685_d N_OUT7_Mp8@1685_g N_VDD_Mp8@1685_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1684 N_OUT8_Mp8@1684_d N_OUT7_Mp8@1684_g N_VDD_Mp8@1684_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1683 N_OUT8_Mn8@1683_d N_OUT7_Mn8@1683_g N_VSS_Mn8@1683_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1682 N_OUT8_Mn8@1682_d N_OUT7_Mn8@1682_g N_VSS_Mn8@1682_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1683 N_OUT8_Mp8@1683_d N_OUT7_Mp8@1683_g N_VDD_Mp8@1683_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1682 N_OUT8_Mp8@1682_d N_OUT7_Mp8@1682_g N_VDD_Mp8@1682_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1681 N_OUT8_Mn8@1681_d N_OUT7_Mn8@1681_g N_VSS_Mn8@1681_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1680 N_OUT8_Mn8@1680_d N_OUT7_Mn8@1680_g N_VSS_Mn8@1680_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1681 N_OUT8_Mp8@1681_d N_OUT7_Mp8@1681_g N_VDD_Mp8@1681_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1680 N_OUT8_Mp8@1680_d N_OUT7_Mp8@1680_g N_VDD_Mp8@1680_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1679 N_OUT8_Mn8@1679_d N_OUT7_Mn8@1679_g N_VSS_Mn8@1679_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1678 N_OUT8_Mn8@1678_d N_OUT7_Mn8@1678_g N_VSS_Mn8@1678_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1679 N_OUT8_Mp8@1679_d N_OUT7_Mp8@1679_g N_VDD_Mp8@1679_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1678 N_OUT8_Mp8@1678_d N_OUT7_Mp8@1678_g N_VDD_Mp8@1678_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1677 N_OUT8_Mn8@1677_d N_OUT7_Mn8@1677_g N_VSS_Mn8@1677_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1676 N_OUT8_Mn8@1676_d N_OUT7_Mn8@1676_g N_VSS_Mn8@1676_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1677 N_OUT8_Mp8@1677_d N_OUT7_Mp8@1677_g N_VDD_Mp8@1677_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1676 N_OUT8_Mp8@1676_d N_OUT7_Mp8@1676_g N_VDD_Mp8@1676_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1675 N_OUT8_Mn8@1675_d N_OUT7_Mn8@1675_g N_VSS_Mn8@1675_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1674 N_OUT8_Mn8@1674_d N_OUT7_Mn8@1674_g N_VSS_Mn8@1674_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1675 N_OUT8_Mp8@1675_d N_OUT7_Mp8@1675_g N_VDD_Mp8@1675_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1674 N_OUT8_Mp8@1674_d N_OUT7_Mp8@1674_g N_VDD_Mp8@1674_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1673 N_OUT8_Mn8@1673_d N_OUT7_Mn8@1673_g N_VSS_Mn8@1673_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1672 N_OUT8_Mn8@1672_d N_OUT7_Mn8@1672_g N_VSS_Mn8@1672_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1673 N_OUT8_Mp8@1673_d N_OUT7_Mp8@1673_g N_VDD_Mp8@1673_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1672 N_OUT8_Mp8@1672_d N_OUT7_Mp8@1672_g N_VDD_Mp8@1672_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1671 N_OUT8_Mn8@1671_d N_OUT7_Mn8@1671_g N_VSS_Mn8@1671_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1670 N_OUT8_Mn8@1670_d N_OUT7_Mn8@1670_g N_VSS_Mn8@1670_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1671 N_OUT8_Mp8@1671_d N_OUT7_Mp8@1671_g N_VDD_Mp8@1671_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1670 N_OUT8_Mp8@1670_d N_OUT7_Mp8@1670_g N_VDD_Mp8@1670_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1669 N_OUT8_Mn8@1669_d N_OUT7_Mn8@1669_g N_VSS_Mn8@1669_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1668 N_OUT8_Mn8@1668_d N_OUT7_Mn8@1668_g N_VSS_Mn8@1668_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1669 N_OUT8_Mp8@1669_d N_OUT7_Mp8@1669_g N_VDD_Mp8@1669_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1668 N_OUT8_Mp8@1668_d N_OUT7_Mp8@1668_g N_VDD_Mp8@1668_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1667 N_OUT8_Mn8@1667_d N_OUT7_Mn8@1667_g N_VSS_Mn8@1667_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1666 N_OUT8_Mn8@1666_d N_OUT7_Mn8@1666_g N_VSS_Mn8@1666_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1667 N_OUT8_Mp8@1667_d N_OUT7_Mp8@1667_g N_VDD_Mp8@1667_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1666 N_OUT8_Mp8@1666_d N_OUT7_Mp8@1666_g N_VDD_Mp8@1666_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1665 N_OUT8_Mn8@1665_d N_OUT7_Mn8@1665_g N_VSS_Mn8@1665_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1664 N_OUT8_Mn8@1664_d N_OUT7_Mn8@1664_g N_VSS_Mn8@1664_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1665 N_OUT8_Mp8@1665_d N_OUT7_Mp8@1665_g N_VDD_Mp8@1665_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1664 N_OUT8_Mp8@1664_d N_OUT7_Mp8@1664_g N_VDD_Mp8@1664_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1663 N_OUT8_Mn8@1663_d N_OUT7_Mn8@1663_g N_VSS_Mn8@1663_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1662 N_OUT8_Mn8@1662_d N_OUT7_Mn8@1662_g N_VSS_Mn8@1662_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1663 N_OUT8_Mp8@1663_d N_OUT7_Mp8@1663_g N_VDD_Mp8@1663_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1662 N_OUT8_Mp8@1662_d N_OUT7_Mp8@1662_g N_VDD_Mp8@1662_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1661 N_OUT8_Mn8@1661_d N_OUT7_Mn8@1661_g N_VSS_Mn8@1661_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1660 N_OUT8_Mn8@1660_d N_OUT7_Mn8@1660_g N_VSS_Mn8@1660_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1661 N_OUT8_Mp8@1661_d N_OUT7_Mp8@1661_g N_VDD_Mp8@1661_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1660 N_OUT8_Mp8@1660_d N_OUT7_Mp8@1660_g N_VDD_Mp8@1660_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1659 N_OUT8_Mn8@1659_d N_OUT7_Mn8@1659_g N_VSS_Mn8@1659_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1658 N_OUT8_Mn8@1658_d N_OUT7_Mn8@1658_g N_VSS_Mn8@1658_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1659 N_OUT8_Mp8@1659_d N_OUT7_Mp8@1659_g N_VDD_Mp8@1659_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1658 N_OUT8_Mp8@1658_d N_OUT7_Mp8@1658_g N_VDD_Mp8@1658_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1657 N_OUT8_Mn8@1657_d N_OUT7_Mn8@1657_g N_VSS_Mn8@1657_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1656 N_OUT8_Mn8@1656_d N_OUT7_Mn8@1656_g N_VSS_Mn8@1656_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1657 N_OUT8_Mp8@1657_d N_OUT7_Mp8@1657_g N_VDD_Mp8@1657_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1656 N_OUT8_Mp8@1656_d N_OUT7_Mp8@1656_g N_VDD_Mp8@1656_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1655 N_OUT8_Mn8@1655_d N_OUT7_Mn8@1655_g N_VSS_Mn8@1655_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1654 N_OUT8_Mn8@1654_d N_OUT7_Mn8@1654_g N_VSS_Mn8@1654_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1655 N_OUT8_Mp8@1655_d N_OUT7_Mp8@1655_g N_VDD_Mp8@1655_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1654 N_OUT8_Mp8@1654_d N_OUT7_Mp8@1654_g N_VDD_Mp8@1654_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1653 N_OUT8_Mn8@1653_d N_OUT7_Mn8@1653_g N_VSS_Mn8@1653_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1652 N_OUT8_Mn8@1652_d N_OUT7_Mn8@1652_g N_VSS_Mn8@1652_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1653 N_OUT8_Mp8@1653_d N_OUT7_Mp8@1653_g N_VDD_Mp8@1653_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1652 N_OUT8_Mp8@1652_d N_OUT7_Mp8@1652_g N_VDD_Mp8@1652_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1651 N_OUT8_Mn8@1651_d N_OUT7_Mn8@1651_g N_VSS_Mn8@1651_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1650 N_OUT8_Mn8@1650_d N_OUT7_Mn8@1650_g N_VSS_Mn8@1650_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1651 N_OUT8_Mp8@1651_d N_OUT7_Mp8@1651_g N_VDD_Mp8@1651_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1650 N_OUT8_Mp8@1650_d N_OUT7_Mp8@1650_g N_VDD_Mp8@1650_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1649 N_OUT8_Mn8@1649_d N_OUT7_Mn8@1649_g N_VSS_Mn8@1649_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1648 N_OUT8_Mn8@1648_d N_OUT7_Mn8@1648_g N_VSS_Mn8@1648_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1649 N_OUT8_Mp8@1649_d N_OUT7_Mp8@1649_g N_VDD_Mp8@1649_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1648 N_OUT8_Mp8@1648_d N_OUT7_Mp8@1648_g N_VDD_Mp8@1648_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1647 N_OUT8_Mn8@1647_d N_OUT7_Mn8@1647_g N_VSS_Mn8@1647_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1646 N_OUT8_Mn8@1646_d N_OUT7_Mn8@1646_g N_VSS_Mn8@1646_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1647 N_OUT8_Mp8@1647_d N_OUT7_Mp8@1647_g N_VDD_Mp8@1647_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1646 N_OUT8_Mp8@1646_d N_OUT7_Mp8@1646_g N_VDD_Mp8@1646_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1645 N_OUT8_Mn8@1645_d N_OUT7_Mn8@1645_g N_VSS_Mn8@1645_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1644 N_OUT8_Mn8@1644_d N_OUT7_Mn8@1644_g N_VSS_Mn8@1644_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1645 N_OUT8_Mp8@1645_d N_OUT7_Mp8@1645_g N_VDD_Mp8@1645_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1644 N_OUT8_Mp8@1644_d N_OUT7_Mp8@1644_g N_VDD_Mp8@1644_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1643 N_OUT8_Mn8@1643_d N_OUT7_Mn8@1643_g N_VSS_Mn8@1643_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1642 N_OUT8_Mn8@1642_d N_OUT7_Mn8@1642_g N_VSS_Mn8@1642_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1643 N_OUT8_Mp8@1643_d N_OUT7_Mp8@1643_g N_VDD_Mp8@1643_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1642 N_OUT8_Mp8@1642_d N_OUT7_Mp8@1642_g N_VDD_Mp8@1642_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1641 N_OUT8_Mn8@1641_d N_OUT7_Mn8@1641_g N_VSS_Mn8@1641_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1640 N_OUT8_Mn8@1640_d N_OUT7_Mn8@1640_g N_VSS_Mn8@1640_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1641 N_OUT8_Mp8@1641_d N_OUT7_Mp8@1641_g N_VDD_Mp8@1641_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1640 N_OUT8_Mp8@1640_d N_OUT7_Mp8@1640_g N_VDD_Mp8@1640_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1639 N_OUT8_Mn8@1639_d N_OUT7_Mn8@1639_g N_VSS_Mn8@1639_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1638 N_OUT8_Mn8@1638_d N_OUT7_Mn8@1638_g N_VSS_Mn8@1638_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1639 N_OUT8_Mp8@1639_d N_OUT7_Mp8@1639_g N_VDD_Mp8@1639_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1638 N_OUT8_Mp8@1638_d N_OUT7_Mp8@1638_g N_VDD_Mp8@1638_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1637 N_OUT8_Mn8@1637_d N_OUT7_Mn8@1637_g N_VSS_Mn8@1637_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1636 N_OUT8_Mn8@1636_d N_OUT7_Mn8@1636_g N_VSS_Mn8@1636_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1637 N_OUT8_Mp8@1637_d N_OUT7_Mp8@1637_g N_VDD_Mp8@1637_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1636 N_OUT8_Mp8@1636_d N_OUT7_Mp8@1636_g N_VDD_Mp8@1636_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1635 N_OUT8_Mn8@1635_d N_OUT7_Mn8@1635_g N_VSS_Mn8@1635_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1634 N_OUT8_Mn8@1634_d N_OUT7_Mn8@1634_g N_VSS_Mn8@1634_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1635 N_OUT8_Mp8@1635_d N_OUT7_Mp8@1635_g N_VDD_Mp8@1635_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1634 N_OUT8_Mp8@1634_d N_OUT7_Mp8@1634_g N_VDD_Mp8@1634_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1633 N_OUT8_Mn8@1633_d N_OUT7_Mn8@1633_g N_VSS_Mn8@1633_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1632 N_OUT8_Mn8@1632_d N_OUT7_Mn8@1632_g N_VSS_Mn8@1632_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1633 N_OUT8_Mp8@1633_d N_OUT7_Mp8@1633_g N_VDD_Mp8@1633_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1632 N_OUT8_Mp8@1632_d N_OUT7_Mp8@1632_g N_VDD_Mp8@1632_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1631 N_OUT8_Mn8@1631_d N_OUT7_Mn8@1631_g N_VSS_Mn8@1631_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1630 N_OUT8_Mn8@1630_d N_OUT7_Mn8@1630_g N_VSS_Mn8@1630_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1631 N_OUT8_Mp8@1631_d N_OUT7_Mp8@1631_g N_VDD_Mp8@1631_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1630 N_OUT8_Mp8@1630_d N_OUT7_Mp8@1630_g N_VDD_Mp8@1630_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1629 N_OUT8_Mn8@1629_d N_OUT7_Mn8@1629_g N_VSS_Mn8@1629_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1628 N_OUT8_Mn8@1628_d N_OUT7_Mn8@1628_g N_VSS_Mn8@1628_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1629 N_OUT8_Mp8@1629_d N_OUT7_Mp8@1629_g N_VDD_Mp8@1629_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1628 N_OUT8_Mp8@1628_d N_OUT7_Mp8@1628_g N_VDD_Mp8@1628_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1627 N_OUT8_Mn8@1627_d N_OUT7_Mn8@1627_g N_VSS_Mn8@1627_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1626 N_OUT8_Mn8@1626_d N_OUT7_Mn8@1626_g N_VSS_Mn8@1626_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1627 N_OUT8_Mp8@1627_d N_OUT7_Mp8@1627_g N_VDD_Mp8@1627_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1626 N_OUT8_Mp8@1626_d N_OUT7_Mp8@1626_g N_VDD_Mp8@1626_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1625 N_OUT8_Mn8@1625_d N_OUT7_Mn8@1625_g N_VSS_Mn8@1625_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1624 N_OUT8_Mn8@1624_d N_OUT7_Mn8@1624_g N_VSS_Mn8@1624_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1625 N_OUT8_Mp8@1625_d N_OUT7_Mp8@1625_g N_VDD_Mp8@1625_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1624 N_OUT8_Mp8@1624_d N_OUT7_Mp8@1624_g N_VDD_Mp8@1624_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1623 N_OUT8_Mn8@1623_d N_OUT7_Mn8@1623_g N_VSS_Mn8@1623_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1622 N_OUT8_Mn8@1622_d N_OUT7_Mn8@1622_g N_VSS_Mn8@1622_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1623 N_OUT8_Mp8@1623_d N_OUT7_Mp8@1623_g N_VDD_Mp8@1623_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1622 N_OUT8_Mp8@1622_d N_OUT7_Mp8@1622_g N_VDD_Mp8@1622_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1621 N_OUT8_Mn8@1621_d N_OUT7_Mn8@1621_g N_VSS_Mn8@1621_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1620 N_OUT8_Mn8@1620_d N_OUT7_Mn8@1620_g N_VSS_Mn8@1620_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1621 N_OUT8_Mp8@1621_d N_OUT7_Mp8@1621_g N_VDD_Mp8@1621_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1620 N_OUT8_Mp8@1620_d N_OUT7_Mp8@1620_g N_VDD_Mp8@1620_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1619 N_OUT8_Mn8@1619_d N_OUT7_Mn8@1619_g N_VSS_Mn8@1619_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1618 N_OUT8_Mn8@1618_d N_OUT7_Mn8@1618_g N_VSS_Mn8@1618_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1619 N_OUT8_Mp8@1619_d N_OUT7_Mp8@1619_g N_VDD_Mp8@1619_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1618 N_OUT8_Mp8@1618_d N_OUT7_Mp8@1618_g N_VDD_Mp8@1618_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1617 N_OUT8_Mn8@1617_d N_OUT7_Mn8@1617_g N_VSS_Mn8@1617_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1616 N_OUT8_Mn8@1616_d N_OUT7_Mn8@1616_g N_VSS_Mn8@1616_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1617 N_OUT8_Mp8@1617_d N_OUT7_Mp8@1617_g N_VDD_Mp8@1617_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1616 N_OUT8_Mp8@1616_d N_OUT7_Mp8@1616_g N_VDD_Mp8@1616_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1615 N_OUT8_Mn8@1615_d N_OUT7_Mn8@1615_g N_VSS_Mn8@1615_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1614 N_OUT8_Mn8@1614_d N_OUT7_Mn8@1614_g N_VSS_Mn8@1614_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1615 N_OUT8_Mp8@1615_d N_OUT7_Mp8@1615_g N_VDD_Mp8@1615_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1614 N_OUT8_Mp8@1614_d N_OUT7_Mp8@1614_g N_VDD_Mp8@1614_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1613 N_OUT8_Mn8@1613_d N_OUT7_Mn8@1613_g N_VSS_Mn8@1613_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1612 N_OUT8_Mn8@1612_d N_OUT7_Mn8@1612_g N_VSS_Mn8@1612_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1613 N_OUT8_Mp8@1613_d N_OUT7_Mp8@1613_g N_VDD_Mp8@1613_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1612 N_OUT8_Mp8@1612_d N_OUT7_Mp8@1612_g N_VDD_Mp8@1612_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1611 N_OUT8_Mn8@1611_d N_OUT7_Mn8@1611_g N_VSS_Mn8@1611_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1610 N_OUT8_Mn8@1610_d N_OUT7_Mn8@1610_g N_VSS_Mn8@1610_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1611 N_OUT8_Mp8@1611_d N_OUT7_Mp8@1611_g N_VDD_Mp8@1611_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1610 N_OUT8_Mp8@1610_d N_OUT7_Mp8@1610_g N_VDD_Mp8@1610_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1609 N_OUT8_Mn8@1609_d N_OUT7_Mn8@1609_g N_VSS_Mn8@1609_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1608 N_OUT8_Mn8@1608_d N_OUT7_Mn8@1608_g N_VSS_Mn8@1608_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1609 N_OUT8_Mp8@1609_d N_OUT7_Mp8@1609_g N_VDD_Mp8@1609_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1608 N_OUT8_Mp8@1608_d N_OUT7_Mp8@1608_g N_VDD_Mp8@1608_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1607 N_OUT8_Mn8@1607_d N_OUT7_Mn8@1607_g N_VSS_Mn8@1607_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1606 N_OUT8_Mn8@1606_d N_OUT7_Mn8@1606_g N_VSS_Mn8@1606_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1607 N_OUT8_Mp8@1607_d N_OUT7_Mp8@1607_g N_VDD_Mp8@1607_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1606 N_OUT8_Mp8@1606_d N_OUT7_Mp8@1606_g N_VDD_Mp8@1606_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1605 N_OUT8_Mn8@1605_d N_OUT7_Mn8@1605_g N_VSS_Mn8@1605_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1604 N_OUT8_Mn8@1604_d N_OUT7_Mn8@1604_g N_VSS_Mn8@1604_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1605 N_OUT8_Mp8@1605_d N_OUT7_Mp8@1605_g N_VDD_Mp8@1605_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1604 N_OUT8_Mp8@1604_d N_OUT7_Mp8@1604_g N_VDD_Mp8@1604_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1603 N_OUT8_Mn8@1603_d N_OUT7_Mn8@1603_g N_VSS_Mn8@1603_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1602 N_OUT8_Mn8@1602_d N_OUT7_Mn8@1602_g N_VSS_Mn8@1602_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1603 N_OUT8_Mp8@1603_d N_OUT7_Mp8@1603_g N_VDD_Mp8@1603_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1602 N_OUT8_Mp8@1602_d N_OUT7_Mp8@1602_g N_VDD_Mp8@1602_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1601 N_OUT8_Mn8@1601_d N_OUT7_Mn8@1601_g N_VSS_Mn8@1601_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1600 N_OUT8_Mn8@1600_d N_OUT7_Mn8@1600_g N_VSS_Mn8@1600_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1601 N_OUT8_Mp8@1601_d N_OUT7_Mp8@1601_g N_VDD_Mp8@1601_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1600 N_OUT8_Mp8@1600_d N_OUT7_Mp8@1600_g N_VDD_Mp8@1600_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1599 N_OUT8_Mn8@1599_d N_OUT7_Mn8@1599_g N_VSS_Mn8@1599_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1598 N_OUT8_Mn8@1598_d N_OUT7_Mn8@1598_g N_VSS_Mn8@1598_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1599 N_OUT8_Mp8@1599_d N_OUT7_Mp8@1599_g N_VDD_Mp8@1599_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1598 N_OUT8_Mp8@1598_d N_OUT7_Mp8@1598_g N_VDD_Mp8@1598_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1597 N_OUT8_Mn8@1597_d N_OUT7_Mn8@1597_g N_VSS_Mn8@1597_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1596 N_OUT8_Mn8@1596_d N_OUT7_Mn8@1596_g N_VSS_Mn8@1596_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1597 N_OUT8_Mp8@1597_d N_OUT7_Mp8@1597_g N_VDD_Mp8@1597_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1596 N_OUT8_Mp8@1596_d N_OUT7_Mp8@1596_g N_VDD_Mp8@1596_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1595 N_OUT8_Mn8@1595_d N_OUT7_Mn8@1595_g N_VSS_Mn8@1595_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1594 N_OUT8_Mn8@1594_d N_OUT7_Mn8@1594_g N_VSS_Mn8@1594_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1595 N_OUT8_Mp8@1595_d N_OUT7_Mp8@1595_g N_VDD_Mp8@1595_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1594 N_OUT8_Mp8@1594_d N_OUT7_Mp8@1594_g N_VDD_Mp8@1594_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1593 N_OUT8_Mn8@1593_d N_OUT7_Mn8@1593_g N_VSS_Mn8@1593_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1592 N_OUT8_Mn8@1592_d N_OUT7_Mn8@1592_g N_VSS_Mn8@1592_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1593 N_OUT8_Mp8@1593_d N_OUT7_Mp8@1593_g N_VDD_Mp8@1593_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1592 N_OUT8_Mp8@1592_d N_OUT7_Mp8@1592_g N_VDD_Mp8@1592_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1591 N_OUT8_Mn8@1591_d N_OUT7_Mn8@1591_g N_VSS_Mn8@1591_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1590 N_OUT8_Mn8@1590_d N_OUT7_Mn8@1590_g N_VSS_Mn8@1590_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1591 N_OUT8_Mp8@1591_d N_OUT7_Mp8@1591_g N_VDD_Mp8@1591_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1590 N_OUT8_Mp8@1590_d N_OUT7_Mp8@1590_g N_VDD_Mp8@1590_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1589 N_OUT8_Mn8@1589_d N_OUT7_Mn8@1589_g N_VSS_Mn8@1589_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1588 N_OUT8_Mn8@1588_d N_OUT7_Mn8@1588_g N_VSS_Mn8@1588_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1589 N_OUT8_Mp8@1589_d N_OUT7_Mp8@1589_g N_VDD_Mp8@1589_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1588 N_OUT8_Mp8@1588_d N_OUT7_Mp8@1588_g N_VDD_Mp8@1588_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1587 N_OUT8_Mn8@1587_d N_OUT7_Mn8@1587_g N_VSS_Mn8@1587_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1586 N_OUT8_Mn8@1586_d N_OUT7_Mn8@1586_g N_VSS_Mn8@1586_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1587 N_OUT8_Mp8@1587_d N_OUT7_Mp8@1587_g N_VDD_Mp8@1587_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1586 N_OUT8_Mp8@1586_d N_OUT7_Mp8@1586_g N_VDD_Mp8@1586_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1585 N_OUT8_Mn8@1585_d N_OUT7_Mn8@1585_g N_VSS_Mn8@1585_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1584 N_OUT8_Mn8@1584_d N_OUT7_Mn8@1584_g N_VSS_Mn8@1584_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1585 N_OUT8_Mp8@1585_d N_OUT7_Mp8@1585_g N_VDD_Mp8@1585_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1584 N_OUT8_Mp8@1584_d N_OUT7_Mp8@1584_g N_VDD_Mp8@1584_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1583 N_OUT8_Mn8@1583_d N_OUT7_Mn8@1583_g N_VSS_Mn8@1583_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1582 N_OUT8_Mn8@1582_d N_OUT7_Mn8@1582_g N_VSS_Mn8@1582_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1583 N_OUT8_Mp8@1583_d N_OUT7_Mp8@1583_g N_VDD_Mp8@1583_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1582 N_OUT8_Mp8@1582_d N_OUT7_Mp8@1582_g N_VDD_Mp8@1582_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1581 N_OUT8_Mn8@1581_d N_OUT7_Mn8@1581_g N_VSS_Mn8@1581_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1580 N_OUT8_Mn8@1580_d N_OUT7_Mn8@1580_g N_VSS_Mn8@1580_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1581 N_OUT8_Mp8@1581_d N_OUT7_Mp8@1581_g N_VDD_Mp8@1581_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1580 N_OUT8_Mp8@1580_d N_OUT7_Mp8@1580_g N_VDD_Mp8@1580_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1579 N_OUT8_Mn8@1579_d N_OUT7_Mn8@1579_g N_VSS_Mn8@1579_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1578 N_OUT8_Mn8@1578_d N_OUT7_Mn8@1578_g N_VSS_Mn8@1578_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1579 N_OUT8_Mp8@1579_d N_OUT7_Mp8@1579_g N_VDD_Mp8@1579_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1578 N_OUT8_Mp8@1578_d N_OUT7_Mp8@1578_g N_VDD_Mp8@1578_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1577 N_OUT8_Mn8@1577_d N_OUT7_Mn8@1577_g N_VSS_Mn8@1577_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1576 N_OUT8_Mn8@1576_d N_OUT7_Mn8@1576_g N_VSS_Mn8@1576_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1577 N_OUT8_Mp8@1577_d N_OUT7_Mp8@1577_g N_VDD_Mp8@1577_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1576 N_OUT8_Mp8@1576_d N_OUT7_Mp8@1576_g N_VDD_Mp8@1576_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1575 N_OUT8_Mn8@1575_d N_OUT7_Mn8@1575_g N_VSS_Mn8@1575_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1574 N_OUT8_Mn8@1574_d N_OUT7_Mn8@1574_g N_VSS_Mn8@1574_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1575 N_OUT8_Mp8@1575_d N_OUT7_Mp8@1575_g N_VDD_Mp8@1575_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1574 N_OUT8_Mp8@1574_d N_OUT7_Mp8@1574_g N_VDD_Mp8@1574_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1573 N_OUT8_Mn8@1573_d N_OUT7_Mn8@1573_g N_VSS_Mn8@1573_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1572 N_OUT8_Mn8@1572_d N_OUT7_Mn8@1572_g N_VSS_Mn8@1572_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1573 N_OUT8_Mp8@1573_d N_OUT7_Mp8@1573_g N_VDD_Mp8@1573_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1572 N_OUT8_Mp8@1572_d N_OUT7_Mp8@1572_g N_VDD_Mp8@1572_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1571 N_OUT8_Mn8@1571_d N_OUT7_Mn8@1571_g N_VSS_Mn8@1571_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1570 N_OUT8_Mn8@1570_d N_OUT7_Mn8@1570_g N_VSS_Mn8@1570_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1571 N_OUT8_Mp8@1571_d N_OUT7_Mp8@1571_g N_VDD_Mp8@1571_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1570 N_OUT8_Mp8@1570_d N_OUT7_Mp8@1570_g N_VDD_Mp8@1570_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1569 N_OUT8_Mn8@1569_d N_OUT7_Mn8@1569_g N_VSS_Mn8@1569_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1568 N_OUT8_Mn8@1568_d N_OUT7_Mn8@1568_g N_VSS_Mn8@1568_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1569 N_OUT8_Mp8@1569_d N_OUT7_Mp8@1569_g N_VDD_Mp8@1569_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1568 N_OUT8_Mp8@1568_d N_OUT7_Mp8@1568_g N_VDD_Mp8@1568_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1567 N_OUT8_Mn8@1567_d N_OUT7_Mn8@1567_g N_VSS_Mn8@1567_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1566 N_OUT8_Mn8@1566_d N_OUT7_Mn8@1566_g N_VSS_Mn8@1566_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1567 N_OUT8_Mp8@1567_d N_OUT7_Mp8@1567_g N_VDD_Mp8@1567_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1566 N_OUT8_Mp8@1566_d N_OUT7_Mp8@1566_g N_VDD_Mp8@1566_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1565 N_OUT8_Mn8@1565_d N_OUT7_Mn8@1565_g N_VSS_Mn8@1565_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1564 N_OUT8_Mn8@1564_d N_OUT7_Mn8@1564_g N_VSS_Mn8@1564_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1565 N_OUT8_Mp8@1565_d N_OUT7_Mp8@1565_g N_VDD_Mp8@1565_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1564 N_OUT8_Mp8@1564_d N_OUT7_Mp8@1564_g N_VDD_Mp8@1564_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1563 N_OUT8_Mn8@1563_d N_OUT7_Mn8@1563_g N_VSS_Mn8@1563_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1562 N_OUT8_Mn8@1562_d N_OUT7_Mn8@1562_g N_VSS_Mn8@1562_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1563 N_OUT8_Mp8@1563_d N_OUT7_Mp8@1563_g N_VDD_Mp8@1563_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1562 N_OUT8_Mp8@1562_d N_OUT7_Mp8@1562_g N_VDD_Mp8@1562_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1561 N_OUT8_Mn8@1561_d N_OUT7_Mn8@1561_g N_VSS_Mn8@1561_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1560 N_OUT8_Mn8@1560_d N_OUT7_Mn8@1560_g N_VSS_Mn8@1560_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1561 N_OUT8_Mp8@1561_d N_OUT7_Mp8@1561_g N_VDD_Mp8@1561_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1560 N_OUT8_Mp8@1560_d N_OUT7_Mp8@1560_g N_VDD_Mp8@1560_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1559 N_OUT8_Mn8@1559_d N_OUT7_Mn8@1559_g N_VSS_Mn8@1559_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1558 N_OUT8_Mn8@1558_d N_OUT7_Mn8@1558_g N_VSS_Mn8@1558_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1559 N_OUT8_Mp8@1559_d N_OUT7_Mp8@1559_g N_VDD_Mp8@1559_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1558 N_OUT8_Mp8@1558_d N_OUT7_Mp8@1558_g N_VDD_Mp8@1558_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1557 N_OUT8_Mn8@1557_d N_OUT7_Mn8@1557_g N_VSS_Mn8@1557_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1556 N_OUT8_Mn8@1556_d N_OUT7_Mn8@1556_g N_VSS_Mn8@1556_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1557 N_OUT8_Mp8@1557_d N_OUT7_Mp8@1557_g N_VDD_Mp8@1557_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1556 N_OUT8_Mp8@1556_d N_OUT7_Mp8@1556_g N_VDD_Mp8@1556_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1555 N_OUT8_Mn8@1555_d N_OUT7_Mn8@1555_g N_VSS_Mn8@1555_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1554 N_OUT8_Mn8@1554_d N_OUT7_Mn8@1554_g N_VSS_Mn8@1554_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1555 N_OUT8_Mp8@1555_d N_OUT7_Mp8@1555_g N_VDD_Mp8@1555_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1554 N_OUT8_Mp8@1554_d N_OUT7_Mp8@1554_g N_VDD_Mp8@1554_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1553 N_OUT8_Mn8@1553_d N_OUT7_Mn8@1553_g N_VSS_Mn8@1553_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1552 N_OUT8_Mn8@1552_d N_OUT7_Mn8@1552_g N_VSS_Mn8@1552_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1553 N_OUT8_Mp8@1553_d N_OUT7_Mp8@1553_g N_VDD_Mp8@1553_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1552 N_OUT8_Mp8@1552_d N_OUT7_Mp8@1552_g N_VDD_Mp8@1552_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1551 N_OUT8_Mn8@1551_d N_OUT7_Mn8@1551_g N_VSS_Mn8@1551_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1550 N_OUT8_Mn8@1550_d N_OUT7_Mn8@1550_g N_VSS_Mn8@1550_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1551 N_OUT8_Mp8@1551_d N_OUT7_Mp8@1551_g N_VDD_Mp8@1551_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1550 N_OUT8_Mp8@1550_d N_OUT7_Mp8@1550_g N_VDD_Mp8@1550_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1549 N_OUT8_Mn8@1549_d N_OUT7_Mn8@1549_g N_VSS_Mn8@1549_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1548 N_OUT8_Mn8@1548_d N_OUT7_Mn8@1548_g N_VSS_Mn8@1548_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1549 N_OUT8_Mp8@1549_d N_OUT7_Mp8@1549_g N_VDD_Mp8@1549_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1548 N_OUT8_Mp8@1548_d N_OUT7_Mp8@1548_g N_VDD_Mp8@1548_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1547 N_OUT8_Mn8@1547_d N_OUT7_Mn8@1547_g N_VSS_Mn8@1547_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1546 N_OUT8_Mn8@1546_d N_OUT7_Mn8@1546_g N_VSS_Mn8@1546_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1547 N_OUT8_Mp8@1547_d N_OUT7_Mp8@1547_g N_VDD_Mp8@1547_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1546 N_OUT8_Mp8@1546_d N_OUT7_Mp8@1546_g N_VDD_Mp8@1546_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1545 N_OUT8_Mn8@1545_d N_OUT7_Mn8@1545_g N_VSS_Mn8@1545_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1544 N_OUT8_Mn8@1544_d N_OUT7_Mn8@1544_g N_VSS_Mn8@1544_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1545 N_OUT8_Mp8@1545_d N_OUT7_Mp8@1545_g N_VDD_Mp8@1545_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1544 N_OUT8_Mp8@1544_d N_OUT7_Mp8@1544_g N_VDD_Mp8@1544_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1543 N_OUT8_Mn8@1543_d N_OUT7_Mn8@1543_g N_VSS_Mn8@1543_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1542 N_OUT8_Mn8@1542_d N_OUT7_Mn8@1542_g N_VSS_Mn8@1542_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1543 N_OUT8_Mp8@1543_d N_OUT7_Mp8@1543_g N_VDD_Mp8@1543_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1542 N_OUT8_Mp8@1542_d N_OUT7_Mp8@1542_g N_VDD_Mp8@1542_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1541 N_OUT8_Mn8@1541_d N_OUT7_Mn8@1541_g N_VSS_Mn8@1541_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1540 N_OUT8_Mn8@1540_d N_OUT7_Mn8@1540_g N_VSS_Mn8@1540_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1541 N_OUT8_Mp8@1541_d N_OUT7_Mp8@1541_g N_VDD_Mp8@1541_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1540 N_OUT8_Mp8@1540_d N_OUT7_Mp8@1540_g N_VDD_Mp8@1540_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1539 N_OUT8_Mn8@1539_d N_OUT7_Mn8@1539_g N_VSS_Mn8@1539_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1538 N_OUT8_Mn8@1538_d N_OUT7_Mn8@1538_g N_VSS_Mn8@1538_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1539 N_OUT8_Mp8@1539_d N_OUT7_Mp8@1539_g N_VDD_Mp8@1539_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1538 N_OUT8_Mp8@1538_d N_OUT7_Mp8@1538_g N_VDD_Mp8@1538_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1537 N_OUT8_Mn8@1537_d N_OUT7_Mn8@1537_g N_VSS_Mn8@1537_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1536 N_OUT8_Mn8@1536_d N_OUT7_Mn8@1536_g N_VSS_Mn8@1536_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1537 N_OUT8_Mp8@1537_d N_OUT7_Mp8@1537_g N_VDD_Mp8@1537_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1536 N_OUT8_Mp8@1536_d N_OUT7_Mp8@1536_g N_VDD_Mp8@1536_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1535 N_OUT8_Mn8@1535_d N_OUT7_Mn8@1535_g N_VSS_Mn8@1535_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1534 N_OUT8_Mn8@1534_d N_OUT7_Mn8@1534_g N_VSS_Mn8@1534_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1535 N_OUT8_Mp8@1535_d N_OUT7_Mp8@1535_g N_VDD_Mp8@1535_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1534 N_OUT8_Mp8@1534_d N_OUT7_Mp8@1534_g N_VDD_Mp8@1534_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1533 N_OUT8_Mn8@1533_d N_OUT7_Mn8@1533_g N_VSS_Mn8@1533_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1532 N_OUT8_Mn8@1532_d N_OUT7_Mn8@1532_g N_VSS_Mn8@1532_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1533 N_OUT8_Mp8@1533_d N_OUT7_Mp8@1533_g N_VDD_Mp8@1533_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1532 N_OUT8_Mp8@1532_d N_OUT7_Mp8@1532_g N_VDD_Mp8@1532_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1531 N_OUT8_Mn8@1531_d N_OUT7_Mn8@1531_g N_VSS_Mn8@1531_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1530 N_OUT8_Mn8@1530_d N_OUT7_Mn8@1530_g N_VSS_Mn8@1530_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1531 N_OUT8_Mp8@1531_d N_OUT7_Mp8@1531_g N_VDD_Mp8@1531_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1530 N_OUT8_Mp8@1530_d N_OUT7_Mp8@1530_g N_VDD_Mp8@1530_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1529 N_OUT8_Mn8@1529_d N_OUT7_Mn8@1529_g N_VSS_Mn8@1529_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1528 N_OUT8_Mn8@1528_d N_OUT7_Mn8@1528_g N_VSS_Mn8@1528_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1529 N_OUT8_Mp8@1529_d N_OUT7_Mp8@1529_g N_VDD_Mp8@1529_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1528 N_OUT8_Mp8@1528_d N_OUT7_Mp8@1528_g N_VDD_Mp8@1528_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1527 N_OUT8_Mn8@1527_d N_OUT7_Mn8@1527_g N_VSS_Mn8@1527_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1526 N_OUT8_Mn8@1526_d N_OUT7_Mn8@1526_g N_VSS_Mn8@1526_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1527 N_OUT8_Mp8@1527_d N_OUT7_Mp8@1527_g N_VDD_Mp8@1527_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1526 N_OUT8_Mp8@1526_d N_OUT7_Mp8@1526_g N_VDD_Mp8@1526_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1525 N_OUT8_Mn8@1525_d N_OUT7_Mn8@1525_g N_VSS_Mn8@1525_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1524 N_OUT8_Mn8@1524_d N_OUT7_Mn8@1524_g N_VSS_Mn8@1524_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1525 N_OUT8_Mp8@1525_d N_OUT7_Mp8@1525_g N_VDD_Mp8@1525_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1524 N_OUT8_Mp8@1524_d N_OUT7_Mp8@1524_g N_VDD_Mp8@1524_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1523 N_OUT8_Mn8@1523_d N_OUT7_Mn8@1523_g N_VSS_Mn8@1523_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1522 N_OUT8_Mn8@1522_d N_OUT7_Mn8@1522_g N_VSS_Mn8@1522_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1523 N_OUT8_Mp8@1523_d N_OUT7_Mp8@1523_g N_VDD_Mp8@1523_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1522 N_OUT8_Mp8@1522_d N_OUT7_Mp8@1522_g N_VDD_Mp8@1522_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1521 N_OUT8_Mn8@1521_d N_OUT7_Mn8@1521_g N_VSS_Mn8@1521_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1520 N_OUT8_Mn8@1520_d N_OUT7_Mn8@1520_g N_VSS_Mn8@1520_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1521 N_OUT8_Mp8@1521_d N_OUT7_Mp8@1521_g N_VDD_Mp8@1521_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1520 N_OUT8_Mp8@1520_d N_OUT7_Mp8@1520_g N_VDD_Mp8@1520_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1519 N_OUT8_Mn8@1519_d N_OUT7_Mn8@1519_g N_VSS_Mn8@1519_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1518 N_OUT8_Mn8@1518_d N_OUT7_Mn8@1518_g N_VSS_Mn8@1518_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1519 N_OUT8_Mp8@1519_d N_OUT7_Mp8@1519_g N_VDD_Mp8@1519_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1518 N_OUT8_Mp8@1518_d N_OUT7_Mp8@1518_g N_VDD_Mp8@1518_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1517 N_OUT8_Mn8@1517_d N_OUT7_Mn8@1517_g N_VSS_Mn8@1517_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1516 N_OUT8_Mn8@1516_d N_OUT7_Mn8@1516_g N_VSS_Mn8@1516_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1517 N_OUT8_Mp8@1517_d N_OUT7_Mp8@1517_g N_VDD_Mp8@1517_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1516 N_OUT8_Mp8@1516_d N_OUT7_Mp8@1516_g N_VDD_Mp8@1516_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1515 N_OUT8_Mn8@1515_d N_OUT7_Mn8@1515_g N_VSS_Mn8@1515_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1514 N_OUT8_Mn8@1514_d N_OUT7_Mn8@1514_g N_VSS_Mn8@1514_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1515 N_OUT8_Mp8@1515_d N_OUT7_Mp8@1515_g N_VDD_Mp8@1515_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1514 N_OUT8_Mp8@1514_d N_OUT7_Mp8@1514_g N_VDD_Mp8@1514_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1513 N_OUT8_Mn8@1513_d N_OUT7_Mn8@1513_g N_VSS_Mn8@1513_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1512 N_OUT8_Mn8@1512_d N_OUT7_Mn8@1512_g N_VSS_Mn8@1512_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1513 N_OUT8_Mp8@1513_d N_OUT7_Mp8@1513_g N_VDD_Mp8@1513_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1512 N_OUT8_Mp8@1512_d N_OUT7_Mp8@1512_g N_VDD_Mp8@1512_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1511 N_OUT8_Mn8@1511_d N_OUT7_Mn8@1511_g N_VSS_Mn8@1511_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1510 N_OUT8_Mn8@1510_d N_OUT7_Mn8@1510_g N_VSS_Mn8@1510_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1511 N_OUT8_Mp8@1511_d N_OUT7_Mp8@1511_g N_VDD_Mp8@1511_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1510 N_OUT8_Mp8@1510_d N_OUT7_Mp8@1510_g N_VDD_Mp8@1510_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1509 N_OUT8_Mn8@1509_d N_OUT7_Mn8@1509_g N_VSS_Mn8@1509_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1508 N_OUT8_Mn8@1508_d N_OUT7_Mn8@1508_g N_VSS_Mn8@1508_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1509 N_OUT8_Mp8@1509_d N_OUT7_Mp8@1509_g N_VDD_Mp8@1509_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1508 N_OUT8_Mp8@1508_d N_OUT7_Mp8@1508_g N_VDD_Mp8@1508_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1507 N_OUT8_Mn8@1507_d N_OUT7_Mn8@1507_g N_VSS_Mn8@1507_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1506 N_OUT8_Mn8@1506_d N_OUT7_Mn8@1506_g N_VSS_Mn8@1506_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1507 N_OUT8_Mp8@1507_d N_OUT7_Mp8@1507_g N_VDD_Mp8@1507_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1506 N_OUT8_Mp8@1506_d N_OUT7_Mp8@1506_g N_VDD_Mp8@1506_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1505 N_OUT8_Mn8@1505_d N_OUT7_Mn8@1505_g N_VSS_Mn8@1505_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1504 N_OUT8_Mn8@1504_d N_OUT7_Mn8@1504_g N_VSS_Mn8@1504_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1505 N_OUT8_Mp8@1505_d N_OUT7_Mp8@1505_g N_VDD_Mp8@1505_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1504 N_OUT8_Mp8@1504_d N_OUT7_Mp8@1504_g N_VDD_Mp8@1504_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1503 N_OUT8_Mn8@1503_d N_OUT7_Mn8@1503_g N_VSS_Mn8@1503_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1502 N_OUT8_Mn8@1502_d N_OUT7_Mn8@1502_g N_VSS_Mn8@1502_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1503 N_OUT8_Mp8@1503_d N_OUT7_Mp8@1503_g N_VDD_Mp8@1503_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1502 N_OUT8_Mp8@1502_d N_OUT7_Mp8@1502_g N_VDD_Mp8@1502_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1501 N_OUT8_Mn8@1501_d N_OUT7_Mn8@1501_g N_VSS_Mn8@1501_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1500 N_OUT8_Mn8@1500_d N_OUT7_Mn8@1500_g N_VSS_Mn8@1500_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1501 N_OUT8_Mp8@1501_d N_OUT7_Mp8@1501_g N_VDD_Mp8@1501_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1500 N_OUT8_Mp8@1500_d N_OUT7_Mp8@1500_g N_VDD_Mp8@1500_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1499 N_OUT8_Mn8@1499_d N_OUT7_Mn8@1499_g N_VSS_Mn8@1499_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1498 N_OUT8_Mn8@1498_d N_OUT7_Mn8@1498_g N_VSS_Mn8@1498_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1499 N_OUT8_Mp8@1499_d N_OUT7_Mp8@1499_g N_VDD_Mp8@1499_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1498 N_OUT8_Mp8@1498_d N_OUT7_Mp8@1498_g N_VDD_Mp8@1498_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1497 N_OUT8_Mn8@1497_d N_OUT7_Mn8@1497_g N_VSS_Mn8@1497_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1496 N_OUT8_Mn8@1496_d N_OUT7_Mn8@1496_g N_VSS_Mn8@1496_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1497 N_OUT8_Mp8@1497_d N_OUT7_Mp8@1497_g N_VDD_Mp8@1497_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1496 N_OUT8_Mp8@1496_d N_OUT7_Mp8@1496_g N_VDD_Mp8@1496_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1495 N_OUT8_Mn8@1495_d N_OUT7_Mn8@1495_g N_VSS_Mn8@1495_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1494 N_OUT8_Mn8@1494_d N_OUT7_Mn8@1494_g N_VSS_Mn8@1494_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1495 N_OUT8_Mp8@1495_d N_OUT7_Mp8@1495_g N_VDD_Mp8@1495_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1494 N_OUT8_Mp8@1494_d N_OUT7_Mp8@1494_g N_VDD_Mp8@1494_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1493 N_OUT8_Mn8@1493_d N_OUT7_Mn8@1493_g N_VSS_Mn8@1493_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1492 N_OUT8_Mn8@1492_d N_OUT7_Mn8@1492_g N_VSS_Mn8@1492_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1493 N_OUT8_Mp8@1493_d N_OUT7_Mp8@1493_g N_VDD_Mp8@1493_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1492 N_OUT8_Mp8@1492_d N_OUT7_Mp8@1492_g N_VDD_Mp8@1492_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1491 N_OUT8_Mn8@1491_d N_OUT7_Mn8@1491_g N_VSS_Mn8@1491_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1490 N_OUT8_Mn8@1490_d N_OUT7_Mn8@1490_g N_VSS_Mn8@1490_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1491 N_OUT8_Mp8@1491_d N_OUT7_Mp8@1491_g N_VDD_Mp8@1491_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1490 N_OUT8_Mp8@1490_d N_OUT7_Mp8@1490_g N_VDD_Mp8@1490_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1489 N_OUT8_Mn8@1489_d N_OUT7_Mn8@1489_g N_VSS_Mn8@1489_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1488 N_OUT8_Mn8@1488_d N_OUT7_Mn8@1488_g N_VSS_Mn8@1488_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1489 N_OUT8_Mp8@1489_d N_OUT7_Mp8@1489_g N_VDD_Mp8@1489_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1488 N_OUT8_Mp8@1488_d N_OUT7_Mp8@1488_g N_VDD_Mp8@1488_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1487 N_OUT8_Mn8@1487_d N_OUT7_Mn8@1487_g N_VSS_Mn8@1487_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1486 N_OUT8_Mn8@1486_d N_OUT7_Mn8@1486_g N_VSS_Mn8@1486_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1487 N_OUT8_Mp8@1487_d N_OUT7_Mp8@1487_g N_VDD_Mp8@1487_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1486 N_OUT8_Mp8@1486_d N_OUT7_Mp8@1486_g N_VDD_Mp8@1486_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1485 N_OUT8_Mn8@1485_d N_OUT7_Mn8@1485_g N_VSS_Mn8@1485_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1484 N_OUT8_Mn8@1484_d N_OUT7_Mn8@1484_g N_VSS_Mn8@1484_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1485 N_OUT8_Mp8@1485_d N_OUT7_Mp8@1485_g N_VDD_Mp8@1485_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1484 N_OUT8_Mp8@1484_d N_OUT7_Mp8@1484_g N_VDD_Mp8@1484_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1483 N_OUT8_Mn8@1483_d N_OUT7_Mn8@1483_g N_VSS_Mn8@1483_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1482 N_OUT8_Mn8@1482_d N_OUT7_Mn8@1482_g N_VSS_Mn8@1482_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1483 N_OUT8_Mp8@1483_d N_OUT7_Mp8@1483_g N_VDD_Mp8@1483_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1482 N_OUT8_Mp8@1482_d N_OUT7_Mp8@1482_g N_VDD_Mp8@1482_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1481 N_OUT8_Mn8@1481_d N_OUT7_Mn8@1481_g N_VSS_Mn8@1481_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1480 N_OUT8_Mn8@1480_d N_OUT7_Mn8@1480_g N_VSS_Mn8@1480_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1481 N_OUT8_Mp8@1481_d N_OUT7_Mp8@1481_g N_VDD_Mp8@1481_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1480 N_OUT8_Mp8@1480_d N_OUT7_Mp8@1480_g N_VDD_Mp8@1480_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1479 N_OUT8_Mn8@1479_d N_OUT7_Mn8@1479_g N_VSS_Mn8@1479_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1478 N_OUT8_Mn8@1478_d N_OUT7_Mn8@1478_g N_VSS_Mn8@1478_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1479 N_OUT8_Mp8@1479_d N_OUT7_Mp8@1479_g N_VDD_Mp8@1479_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1478 N_OUT8_Mp8@1478_d N_OUT7_Mp8@1478_g N_VDD_Mp8@1478_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1477 N_OUT8_Mn8@1477_d N_OUT7_Mn8@1477_g N_VSS_Mn8@1477_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1476 N_OUT8_Mn8@1476_d N_OUT7_Mn8@1476_g N_VSS_Mn8@1476_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1477 N_OUT8_Mp8@1477_d N_OUT7_Mp8@1477_g N_VDD_Mp8@1477_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1476 N_OUT8_Mp8@1476_d N_OUT7_Mp8@1476_g N_VDD_Mp8@1476_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1475 N_OUT8_Mn8@1475_d N_OUT7_Mn8@1475_g N_VSS_Mn8@1475_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1474 N_OUT8_Mn8@1474_d N_OUT7_Mn8@1474_g N_VSS_Mn8@1474_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1475 N_OUT8_Mp8@1475_d N_OUT7_Mp8@1475_g N_VDD_Mp8@1475_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1474 N_OUT8_Mp8@1474_d N_OUT7_Mp8@1474_g N_VDD_Mp8@1474_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1473 N_OUT8_Mn8@1473_d N_OUT7_Mn8@1473_g N_VSS_Mn8@1473_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1472 N_OUT8_Mn8@1472_d N_OUT7_Mn8@1472_g N_VSS_Mn8@1472_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1473 N_OUT8_Mp8@1473_d N_OUT7_Mp8@1473_g N_VDD_Mp8@1473_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1472 N_OUT8_Mp8@1472_d N_OUT7_Mp8@1472_g N_VDD_Mp8@1472_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1471 N_OUT8_Mn8@1471_d N_OUT7_Mn8@1471_g N_VSS_Mn8@1471_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1470 N_OUT8_Mn8@1470_d N_OUT7_Mn8@1470_g N_VSS_Mn8@1470_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1471 N_OUT8_Mp8@1471_d N_OUT7_Mp8@1471_g N_VDD_Mp8@1471_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1470 N_OUT8_Mp8@1470_d N_OUT7_Mp8@1470_g N_VDD_Mp8@1470_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1469 N_OUT8_Mn8@1469_d N_OUT7_Mn8@1469_g N_VSS_Mn8@1469_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1468 N_OUT8_Mn8@1468_d N_OUT7_Mn8@1468_g N_VSS_Mn8@1468_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1469 N_OUT8_Mp8@1469_d N_OUT7_Mp8@1469_g N_VDD_Mp8@1469_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1468 N_OUT8_Mp8@1468_d N_OUT7_Mp8@1468_g N_VDD_Mp8@1468_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1467 N_OUT8_Mn8@1467_d N_OUT7_Mn8@1467_g N_VSS_Mn8@1467_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1466 N_OUT8_Mn8@1466_d N_OUT7_Mn8@1466_g N_VSS_Mn8@1466_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1467 N_OUT8_Mp8@1467_d N_OUT7_Mp8@1467_g N_VDD_Mp8@1467_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1466 N_OUT8_Mp8@1466_d N_OUT7_Mp8@1466_g N_VDD_Mp8@1466_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1465 N_OUT8_Mn8@1465_d N_OUT7_Mn8@1465_g N_VSS_Mn8@1465_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1464 N_OUT8_Mn8@1464_d N_OUT7_Mn8@1464_g N_VSS_Mn8@1464_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1465 N_OUT8_Mp8@1465_d N_OUT7_Mp8@1465_g N_VDD_Mp8@1465_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1464 N_OUT8_Mp8@1464_d N_OUT7_Mp8@1464_g N_VDD_Mp8@1464_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1463 N_OUT8_Mn8@1463_d N_OUT7_Mn8@1463_g N_VSS_Mn8@1463_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1462 N_OUT8_Mn8@1462_d N_OUT7_Mn8@1462_g N_VSS_Mn8@1462_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1463 N_OUT8_Mp8@1463_d N_OUT7_Mp8@1463_g N_VDD_Mp8@1463_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1462 N_OUT8_Mp8@1462_d N_OUT7_Mp8@1462_g N_VDD_Mp8@1462_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1461 N_OUT8_Mn8@1461_d N_OUT7_Mn8@1461_g N_VSS_Mn8@1461_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1460 N_OUT8_Mn8@1460_d N_OUT7_Mn8@1460_g N_VSS_Mn8@1460_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1461 N_OUT8_Mp8@1461_d N_OUT7_Mp8@1461_g N_VDD_Mp8@1461_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1460 N_OUT8_Mp8@1460_d N_OUT7_Mp8@1460_g N_VDD_Mp8@1460_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1459 N_OUT8_Mn8@1459_d N_OUT7_Mn8@1459_g N_VSS_Mn8@1459_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1458 N_OUT8_Mn8@1458_d N_OUT7_Mn8@1458_g N_VSS_Mn8@1458_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1459 N_OUT8_Mp8@1459_d N_OUT7_Mp8@1459_g N_VDD_Mp8@1459_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1458 N_OUT8_Mp8@1458_d N_OUT7_Mp8@1458_g N_VDD_Mp8@1458_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1457 N_OUT8_Mn8@1457_d N_OUT7_Mn8@1457_g N_VSS_Mn8@1457_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1456 N_OUT8_Mn8@1456_d N_OUT7_Mn8@1456_g N_VSS_Mn8@1456_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1457 N_OUT8_Mp8@1457_d N_OUT7_Mp8@1457_g N_VDD_Mp8@1457_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1456 N_OUT8_Mp8@1456_d N_OUT7_Mp8@1456_g N_VDD_Mp8@1456_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1455 N_OUT8_Mn8@1455_d N_OUT7_Mn8@1455_g N_VSS_Mn8@1455_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1454 N_OUT8_Mn8@1454_d N_OUT7_Mn8@1454_g N_VSS_Mn8@1454_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1455 N_OUT8_Mp8@1455_d N_OUT7_Mp8@1455_g N_VDD_Mp8@1455_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1454 N_OUT8_Mp8@1454_d N_OUT7_Mp8@1454_g N_VDD_Mp8@1454_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1453 N_OUT8_Mn8@1453_d N_OUT7_Mn8@1453_g N_VSS_Mn8@1453_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1452 N_OUT8_Mn8@1452_d N_OUT7_Mn8@1452_g N_VSS_Mn8@1452_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1453 N_OUT8_Mp8@1453_d N_OUT7_Mp8@1453_g N_VDD_Mp8@1453_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1452 N_OUT8_Mp8@1452_d N_OUT7_Mp8@1452_g N_VDD_Mp8@1452_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1451 N_OUT8_Mn8@1451_d N_OUT7_Mn8@1451_g N_VSS_Mn8@1451_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1450 N_OUT8_Mn8@1450_d N_OUT7_Mn8@1450_g N_VSS_Mn8@1450_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1451 N_OUT8_Mp8@1451_d N_OUT7_Mp8@1451_g N_VDD_Mp8@1451_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1450 N_OUT8_Mp8@1450_d N_OUT7_Mp8@1450_g N_VDD_Mp8@1450_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1449 N_OUT8_Mn8@1449_d N_OUT7_Mn8@1449_g N_VSS_Mn8@1449_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1448 N_OUT8_Mn8@1448_d N_OUT7_Mn8@1448_g N_VSS_Mn8@1448_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1449 N_OUT8_Mp8@1449_d N_OUT7_Mp8@1449_g N_VDD_Mp8@1449_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1448 N_OUT8_Mp8@1448_d N_OUT7_Mp8@1448_g N_VDD_Mp8@1448_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1447 N_OUT8_Mn8@1447_d N_OUT7_Mn8@1447_g N_VSS_Mn8@1447_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1446 N_OUT8_Mn8@1446_d N_OUT7_Mn8@1446_g N_VSS_Mn8@1446_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1447 N_OUT8_Mp8@1447_d N_OUT7_Mp8@1447_g N_VDD_Mp8@1447_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1446 N_OUT8_Mp8@1446_d N_OUT7_Mp8@1446_g N_VDD_Mp8@1446_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1445 N_OUT8_Mn8@1445_d N_OUT7_Mn8@1445_g N_VSS_Mn8@1445_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1444 N_OUT8_Mn8@1444_d N_OUT7_Mn8@1444_g N_VSS_Mn8@1444_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1445 N_OUT8_Mp8@1445_d N_OUT7_Mp8@1445_g N_VDD_Mp8@1445_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1444 N_OUT8_Mp8@1444_d N_OUT7_Mp8@1444_g N_VDD_Mp8@1444_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1443 N_OUT8_Mn8@1443_d N_OUT7_Mn8@1443_g N_VSS_Mn8@1443_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1442 N_OUT8_Mn8@1442_d N_OUT7_Mn8@1442_g N_VSS_Mn8@1442_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1443 N_OUT8_Mp8@1443_d N_OUT7_Mp8@1443_g N_VDD_Mp8@1443_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1442 N_OUT8_Mp8@1442_d N_OUT7_Mp8@1442_g N_VDD_Mp8@1442_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1441 N_OUT8_Mn8@1441_d N_OUT7_Mn8@1441_g N_VSS_Mn8@1441_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1440 N_OUT8_Mn8@1440_d N_OUT7_Mn8@1440_g N_VSS_Mn8@1440_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1441 N_OUT8_Mp8@1441_d N_OUT7_Mp8@1441_g N_VDD_Mp8@1441_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1440 N_OUT8_Mp8@1440_d N_OUT7_Mp8@1440_g N_VDD_Mp8@1440_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1439 N_OUT8_Mn8@1439_d N_OUT7_Mn8@1439_g N_VSS_Mn8@1439_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1438 N_OUT8_Mn8@1438_d N_OUT7_Mn8@1438_g N_VSS_Mn8@1438_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1439 N_OUT8_Mp8@1439_d N_OUT7_Mp8@1439_g N_VDD_Mp8@1439_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1438 N_OUT8_Mp8@1438_d N_OUT7_Mp8@1438_g N_VDD_Mp8@1438_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1437 N_OUT8_Mn8@1437_d N_OUT7_Mn8@1437_g N_VSS_Mn8@1437_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1436 N_OUT8_Mn8@1436_d N_OUT7_Mn8@1436_g N_VSS_Mn8@1436_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1437 N_OUT8_Mp8@1437_d N_OUT7_Mp8@1437_g N_VDD_Mp8@1437_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1436 N_OUT8_Mp8@1436_d N_OUT7_Mp8@1436_g N_VDD_Mp8@1436_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1435 N_OUT8_Mn8@1435_d N_OUT7_Mn8@1435_g N_VSS_Mn8@1435_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1434 N_OUT8_Mn8@1434_d N_OUT7_Mn8@1434_g N_VSS_Mn8@1434_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1435 N_OUT8_Mp8@1435_d N_OUT7_Mp8@1435_g N_VDD_Mp8@1435_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1434 N_OUT8_Mp8@1434_d N_OUT7_Mp8@1434_g N_VDD_Mp8@1434_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1433 N_OUT8_Mn8@1433_d N_OUT7_Mn8@1433_g N_VSS_Mn8@1433_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1432 N_OUT8_Mn8@1432_d N_OUT7_Mn8@1432_g N_VSS_Mn8@1432_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1433 N_OUT8_Mp8@1433_d N_OUT7_Mp8@1433_g N_VDD_Mp8@1433_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1432 N_OUT8_Mp8@1432_d N_OUT7_Mp8@1432_g N_VDD_Mp8@1432_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1431 N_OUT8_Mn8@1431_d N_OUT7_Mn8@1431_g N_VSS_Mn8@1431_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1430 N_OUT8_Mn8@1430_d N_OUT7_Mn8@1430_g N_VSS_Mn8@1430_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1431 N_OUT8_Mp8@1431_d N_OUT7_Mp8@1431_g N_VDD_Mp8@1431_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1430 N_OUT8_Mp8@1430_d N_OUT7_Mp8@1430_g N_VDD_Mp8@1430_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1429 N_OUT8_Mn8@1429_d N_OUT7_Mn8@1429_g N_VSS_Mn8@1429_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1428 N_OUT8_Mn8@1428_d N_OUT7_Mn8@1428_g N_VSS_Mn8@1428_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1429 N_OUT8_Mp8@1429_d N_OUT7_Mp8@1429_g N_VDD_Mp8@1429_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1428 N_OUT8_Mp8@1428_d N_OUT7_Mp8@1428_g N_VDD_Mp8@1428_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1427 N_OUT8_Mn8@1427_d N_OUT7_Mn8@1427_g N_VSS_Mn8@1427_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1426 N_OUT8_Mn8@1426_d N_OUT7_Mn8@1426_g N_VSS_Mn8@1426_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1427 N_OUT8_Mp8@1427_d N_OUT7_Mp8@1427_g N_VDD_Mp8@1427_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1426 N_OUT8_Mp8@1426_d N_OUT7_Mp8@1426_g N_VDD_Mp8@1426_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1425 N_OUT8_Mn8@1425_d N_OUT7_Mn8@1425_g N_VSS_Mn8@1425_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1424 N_OUT8_Mn8@1424_d N_OUT7_Mn8@1424_g N_VSS_Mn8@1424_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1425 N_OUT8_Mp8@1425_d N_OUT7_Mp8@1425_g N_VDD_Mp8@1425_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1424 N_OUT8_Mp8@1424_d N_OUT7_Mp8@1424_g N_VDD_Mp8@1424_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1423 N_OUT8_Mn8@1423_d N_OUT7_Mn8@1423_g N_VSS_Mn8@1423_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1422 N_OUT8_Mn8@1422_d N_OUT7_Mn8@1422_g N_VSS_Mn8@1422_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1423 N_OUT8_Mp8@1423_d N_OUT7_Mp8@1423_g N_VDD_Mp8@1423_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1422 N_OUT8_Mp8@1422_d N_OUT7_Mp8@1422_g N_VDD_Mp8@1422_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1421 N_OUT8_Mn8@1421_d N_OUT7_Mn8@1421_g N_VSS_Mn8@1421_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1420 N_OUT8_Mn8@1420_d N_OUT7_Mn8@1420_g N_VSS_Mn8@1420_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1421 N_OUT8_Mp8@1421_d N_OUT7_Mp8@1421_g N_VDD_Mp8@1421_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1420 N_OUT8_Mp8@1420_d N_OUT7_Mp8@1420_g N_VDD_Mp8@1420_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1419 N_OUT8_Mn8@1419_d N_OUT7_Mn8@1419_g N_VSS_Mn8@1419_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1418 N_OUT8_Mn8@1418_d N_OUT7_Mn8@1418_g N_VSS_Mn8@1418_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1419 N_OUT8_Mp8@1419_d N_OUT7_Mp8@1419_g N_VDD_Mp8@1419_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1418 N_OUT8_Mp8@1418_d N_OUT7_Mp8@1418_g N_VDD_Mp8@1418_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1417 N_OUT8_Mn8@1417_d N_OUT7_Mn8@1417_g N_VSS_Mn8@1417_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1416 N_OUT8_Mn8@1416_d N_OUT7_Mn8@1416_g N_VSS_Mn8@1416_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1417 N_OUT8_Mp8@1417_d N_OUT7_Mp8@1417_g N_VDD_Mp8@1417_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1416 N_OUT8_Mp8@1416_d N_OUT7_Mp8@1416_g N_VDD_Mp8@1416_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1415 N_OUT8_Mn8@1415_d N_OUT7_Mn8@1415_g N_VSS_Mn8@1415_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1414 N_OUT8_Mn8@1414_d N_OUT7_Mn8@1414_g N_VSS_Mn8@1414_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1415 N_OUT8_Mp8@1415_d N_OUT7_Mp8@1415_g N_VDD_Mp8@1415_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1414 N_OUT8_Mp8@1414_d N_OUT7_Mp8@1414_g N_VDD_Mp8@1414_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1413 N_OUT8_Mn8@1413_d N_OUT7_Mn8@1413_g N_VSS_Mn8@1413_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1412 N_OUT8_Mn8@1412_d N_OUT7_Mn8@1412_g N_VSS_Mn8@1412_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1413 N_OUT8_Mp8@1413_d N_OUT7_Mp8@1413_g N_VDD_Mp8@1413_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1412 N_OUT8_Mp8@1412_d N_OUT7_Mp8@1412_g N_VDD_Mp8@1412_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1411 N_OUT8_Mn8@1411_d N_OUT7_Mn8@1411_g N_VSS_Mn8@1411_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1410 N_OUT8_Mn8@1410_d N_OUT7_Mn8@1410_g N_VSS_Mn8@1410_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1411 N_OUT8_Mp8@1411_d N_OUT7_Mp8@1411_g N_VDD_Mp8@1411_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1410 N_OUT8_Mp8@1410_d N_OUT7_Mp8@1410_g N_VDD_Mp8@1410_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1409 N_OUT8_Mn8@1409_d N_OUT7_Mn8@1409_g N_VSS_Mn8@1409_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1408 N_OUT8_Mn8@1408_d N_OUT7_Mn8@1408_g N_VSS_Mn8@1408_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1409 N_OUT8_Mp8@1409_d N_OUT7_Mp8@1409_g N_VDD_Mp8@1409_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1408 N_OUT8_Mp8@1408_d N_OUT7_Mp8@1408_g N_VDD_Mp8@1408_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1407 N_OUT8_Mn8@1407_d N_OUT7_Mn8@1407_g N_VSS_Mn8@1407_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1406 N_OUT8_Mn8@1406_d N_OUT7_Mn8@1406_g N_VSS_Mn8@1406_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1407 N_OUT8_Mp8@1407_d N_OUT7_Mp8@1407_g N_VDD_Mp8@1407_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1406 N_OUT8_Mp8@1406_d N_OUT7_Mp8@1406_g N_VDD_Mp8@1406_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1405 N_OUT8_Mn8@1405_d N_OUT7_Mn8@1405_g N_VSS_Mn8@1405_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1404 N_OUT8_Mn8@1404_d N_OUT7_Mn8@1404_g N_VSS_Mn8@1404_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1405 N_OUT8_Mp8@1405_d N_OUT7_Mp8@1405_g N_VDD_Mp8@1405_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1404 N_OUT8_Mp8@1404_d N_OUT7_Mp8@1404_g N_VDD_Mp8@1404_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1403 N_OUT8_Mn8@1403_d N_OUT7_Mn8@1403_g N_VSS_Mn8@1403_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1402 N_OUT8_Mn8@1402_d N_OUT7_Mn8@1402_g N_VSS_Mn8@1402_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1403 N_OUT8_Mp8@1403_d N_OUT7_Mp8@1403_g N_VDD_Mp8@1403_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1402 N_OUT8_Mp8@1402_d N_OUT7_Mp8@1402_g N_VDD_Mp8@1402_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1401 N_OUT8_Mn8@1401_d N_OUT7_Mn8@1401_g N_VSS_Mn8@1401_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1400 N_OUT8_Mn8@1400_d N_OUT7_Mn8@1400_g N_VSS_Mn8@1400_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1401 N_OUT8_Mp8@1401_d N_OUT7_Mp8@1401_g N_VDD_Mp8@1401_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1400 N_OUT8_Mp8@1400_d N_OUT7_Mp8@1400_g N_VDD_Mp8@1400_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1399 N_OUT8_Mn8@1399_d N_OUT7_Mn8@1399_g N_VSS_Mn8@1399_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1398 N_OUT8_Mn8@1398_d N_OUT7_Mn8@1398_g N_VSS_Mn8@1398_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1399 N_OUT8_Mp8@1399_d N_OUT7_Mp8@1399_g N_VDD_Mp8@1399_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1398 N_OUT8_Mp8@1398_d N_OUT7_Mp8@1398_g N_VDD_Mp8@1398_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1397 N_OUT8_Mn8@1397_d N_OUT7_Mn8@1397_g N_VSS_Mn8@1397_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1396 N_OUT8_Mn8@1396_d N_OUT7_Mn8@1396_g N_VSS_Mn8@1396_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1397 N_OUT8_Mp8@1397_d N_OUT7_Mp8@1397_g N_VDD_Mp8@1397_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1396 N_OUT8_Mp8@1396_d N_OUT7_Mp8@1396_g N_VDD_Mp8@1396_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1395 N_OUT8_Mn8@1395_d N_OUT7_Mn8@1395_g N_VSS_Mn8@1395_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1394 N_OUT8_Mn8@1394_d N_OUT7_Mn8@1394_g N_VSS_Mn8@1394_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1395 N_OUT8_Mp8@1395_d N_OUT7_Mp8@1395_g N_VDD_Mp8@1395_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1394 N_OUT8_Mp8@1394_d N_OUT7_Mp8@1394_g N_VDD_Mp8@1394_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1393 N_OUT8_Mn8@1393_d N_OUT7_Mn8@1393_g N_VSS_Mn8@1393_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1392 N_OUT8_Mn8@1392_d N_OUT7_Mn8@1392_g N_VSS_Mn8@1392_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1393 N_OUT8_Mp8@1393_d N_OUT7_Mp8@1393_g N_VDD_Mp8@1393_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1392 N_OUT8_Mp8@1392_d N_OUT7_Mp8@1392_g N_VDD_Mp8@1392_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1391 N_OUT8_Mn8@1391_d N_OUT7_Mn8@1391_g N_VSS_Mn8@1391_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1390 N_OUT8_Mn8@1390_d N_OUT7_Mn8@1390_g N_VSS_Mn8@1390_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1391 N_OUT8_Mp8@1391_d N_OUT7_Mp8@1391_g N_VDD_Mp8@1391_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1390 N_OUT8_Mp8@1390_d N_OUT7_Mp8@1390_g N_VDD_Mp8@1390_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1389 N_OUT8_Mn8@1389_d N_OUT7_Mn8@1389_g N_VSS_Mn8@1389_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1388 N_OUT8_Mn8@1388_d N_OUT7_Mn8@1388_g N_VSS_Mn8@1388_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1389 N_OUT8_Mp8@1389_d N_OUT7_Mp8@1389_g N_VDD_Mp8@1389_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1388 N_OUT8_Mp8@1388_d N_OUT7_Mp8@1388_g N_VDD_Mp8@1388_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1387 N_OUT8_Mn8@1387_d N_OUT7_Mn8@1387_g N_VSS_Mn8@1387_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1386 N_OUT8_Mn8@1386_d N_OUT7_Mn8@1386_g N_VSS_Mn8@1386_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1387 N_OUT8_Mp8@1387_d N_OUT7_Mp8@1387_g N_VDD_Mp8@1387_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1386 N_OUT8_Mp8@1386_d N_OUT7_Mp8@1386_g N_VDD_Mp8@1386_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1385 N_OUT8_Mn8@1385_d N_OUT7_Mn8@1385_g N_VSS_Mn8@1385_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1384 N_OUT8_Mn8@1384_d N_OUT7_Mn8@1384_g N_VSS_Mn8@1384_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1385 N_OUT8_Mp8@1385_d N_OUT7_Mp8@1385_g N_VDD_Mp8@1385_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1384 N_OUT8_Mp8@1384_d N_OUT7_Mp8@1384_g N_VDD_Mp8@1384_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1383 N_OUT8_Mn8@1383_d N_OUT7_Mn8@1383_g N_VSS_Mn8@1383_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1382 N_OUT8_Mn8@1382_d N_OUT7_Mn8@1382_g N_VSS_Mn8@1382_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1383 N_OUT8_Mp8@1383_d N_OUT7_Mp8@1383_g N_VDD_Mp8@1383_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1382 N_OUT8_Mp8@1382_d N_OUT7_Mp8@1382_g N_VDD_Mp8@1382_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1381 N_OUT8_Mn8@1381_d N_OUT7_Mn8@1381_g N_VSS_Mn8@1381_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1380 N_OUT8_Mn8@1380_d N_OUT7_Mn8@1380_g N_VSS_Mn8@1380_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1381 N_OUT8_Mp8@1381_d N_OUT7_Mp8@1381_g N_VDD_Mp8@1381_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1380 N_OUT8_Mp8@1380_d N_OUT7_Mp8@1380_g N_VDD_Mp8@1380_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1379 N_OUT8_Mn8@1379_d N_OUT7_Mn8@1379_g N_VSS_Mn8@1379_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1378 N_OUT8_Mn8@1378_d N_OUT7_Mn8@1378_g N_VSS_Mn8@1378_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1379 N_OUT8_Mp8@1379_d N_OUT7_Mp8@1379_g N_VDD_Mp8@1379_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1378 N_OUT8_Mp8@1378_d N_OUT7_Mp8@1378_g N_VDD_Mp8@1378_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1377 N_OUT8_Mn8@1377_d N_OUT7_Mn8@1377_g N_VSS_Mn8@1377_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1376 N_OUT8_Mn8@1376_d N_OUT7_Mn8@1376_g N_VSS_Mn8@1376_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1377 N_OUT8_Mp8@1377_d N_OUT7_Mp8@1377_g N_VDD_Mp8@1377_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1376 N_OUT8_Mp8@1376_d N_OUT7_Mp8@1376_g N_VDD_Mp8@1376_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1375 N_OUT8_Mn8@1375_d N_OUT7_Mn8@1375_g N_VSS_Mn8@1375_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1374 N_OUT8_Mn8@1374_d N_OUT7_Mn8@1374_g N_VSS_Mn8@1374_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1375 N_OUT8_Mp8@1375_d N_OUT7_Mp8@1375_g N_VDD_Mp8@1375_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1374 N_OUT8_Mp8@1374_d N_OUT7_Mp8@1374_g N_VDD_Mp8@1374_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1373 N_OUT8_Mn8@1373_d N_OUT7_Mn8@1373_g N_VSS_Mn8@1373_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1372 N_OUT8_Mn8@1372_d N_OUT7_Mn8@1372_g N_VSS_Mn8@1372_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1373 N_OUT8_Mp8@1373_d N_OUT7_Mp8@1373_g N_VDD_Mp8@1373_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1372 N_OUT8_Mp8@1372_d N_OUT7_Mp8@1372_g N_VDD_Mp8@1372_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1371 N_OUT8_Mn8@1371_d N_OUT7_Mn8@1371_g N_VSS_Mn8@1371_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1370 N_OUT8_Mn8@1370_d N_OUT7_Mn8@1370_g N_VSS_Mn8@1370_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1371 N_OUT8_Mp8@1371_d N_OUT7_Mp8@1371_g N_VDD_Mp8@1371_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1370 N_OUT8_Mp8@1370_d N_OUT7_Mp8@1370_g N_VDD_Mp8@1370_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1369 N_OUT8_Mn8@1369_d N_OUT7_Mn8@1369_g N_VSS_Mn8@1369_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1368 N_OUT8_Mn8@1368_d N_OUT7_Mn8@1368_g N_VSS_Mn8@1368_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1369 N_OUT8_Mp8@1369_d N_OUT7_Mp8@1369_g N_VDD_Mp8@1369_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1368 N_OUT8_Mp8@1368_d N_OUT7_Mp8@1368_g N_VDD_Mp8@1368_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1367 N_OUT8_Mn8@1367_d N_OUT7_Mn8@1367_g N_VSS_Mn8@1367_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1366 N_OUT8_Mn8@1366_d N_OUT7_Mn8@1366_g N_VSS_Mn8@1366_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1367 N_OUT8_Mp8@1367_d N_OUT7_Mp8@1367_g N_VDD_Mp8@1367_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1366 N_OUT8_Mp8@1366_d N_OUT7_Mp8@1366_g N_VDD_Mp8@1366_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1365 N_OUT8_Mn8@1365_d N_OUT7_Mn8@1365_g N_VSS_Mn8@1365_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1364 N_OUT8_Mn8@1364_d N_OUT7_Mn8@1364_g N_VSS_Mn8@1364_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1365 N_OUT8_Mp8@1365_d N_OUT7_Mp8@1365_g N_VDD_Mp8@1365_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1364 N_OUT8_Mp8@1364_d N_OUT7_Mp8@1364_g N_VDD_Mp8@1364_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1363 N_OUT8_Mn8@1363_d N_OUT7_Mn8@1363_g N_VSS_Mn8@1363_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1362 N_OUT8_Mn8@1362_d N_OUT7_Mn8@1362_g N_VSS_Mn8@1362_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1363 N_OUT8_Mp8@1363_d N_OUT7_Mp8@1363_g N_VDD_Mp8@1363_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1362 N_OUT8_Mp8@1362_d N_OUT7_Mp8@1362_g N_VDD_Mp8@1362_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1361 N_OUT8_Mn8@1361_d N_OUT7_Mn8@1361_g N_VSS_Mn8@1361_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1360 N_OUT8_Mn8@1360_d N_OUT7_Mn8@1360_g N_VSS_Mn8@1360_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1361 N_OUT8_Mp8@1361_d N_OUT7_Mp8@1361_g N_VDD_Mp8@1361_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1360 N_OUT8_Mp8@1360_d N_OUT7_Mp8@1360_g N_VDD_Mp8@1360_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1359 N_OUT8_Mn8@1359_d N_OUT7_Mn8@1359_g N_VSS_Mn8@1359_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1358 N_OUT8_Mn8@1358_d N_OUT7_Mn8@1358_g N_VSS_Mn8@1358_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1359 N_OUT8_Mp8@1359_d N_OUT7_Mp8@1359_g N_VDD_Mp8@1359_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1358 N_OUT8_Mp8@1358_d N_OUT7_Mp8@1358_g N_VDD_Mp8@1358_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1357 N_OUT8_Mn8@1357_d N_OUT7_Mn8@1357_g N_VSS_Mn8@1357_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1356 N_OUT8_Mn8@1356_d N_OUT7_Mn8@1356_g N_VSS_Mn8@1356_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1357 N_OUT8_Mp8@1357_d N_OUT7_Mp8@1357_g N_VDD_Mp8@1357_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1356 N_OUT8_Mp8@1356_d N_OUT7_Mp8@1356_g N_VDD_Mp8@1356_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1355 N_OUT8_Mn8@1355_d N_OUT7_Mn8@1355_g N_VSS_Mn8@1355_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1354 N_OUT8_Mn8@1354_d N_OUT7_Mn8@1354_g N_VSS_Mn8@1354_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1355 N_OUT8_Mp8@1355_d N_OUT7_Mp8@1355_g N_VDD_Mp8@1355_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1354 N_OUT8_Mp8@1354_d N_OUT7_Mp8@1354_g N_VDD_Mp8@1354_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1353 N_OUT8_Mn8@1353_d N_OUT7_Mn8@1353_g N_VSS_Mn8@1353_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1352 N_OUT8_Mn8@1352_d N_OUT7_Mn8@1352_g N_VSS_Mn8@1352_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1353 N_OUT8_Mp8@1353_d N_OUT7_Mp8@1353_g N_VDD_Mp8@1353_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1352 N_OUT8_Mp8@1352_d N_OUT7_Mp8@1352_g N_VDD_Mp8@1352_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1351 N_OUT8_Mn8@1351_d N_OUT7_Mn8@1351_g N_VSS_Mn8@1351_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1350 N_OUT8_Mn8@1350_d N_OUT7_Mn8@1350_g N_VSS_Mn8@1350_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1351 N_OUT8_Mp8@1351_d N_OUT7_Mp8@1351_g N_VDD_Mp8@1351_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1350 N_OUT8_Mp8@1350_d N_OUT7_Mp8@1350_g N_VDD_Mp8@1350_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1349 N_OUT8_Mn8@1349_d N_OUT7_Mn8@1349_g N_VSS_Mn8@1349_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1348 N_OUT8_Mn8@1348_d N_OUT7_Mn8@1348_g N_VSS_Mn8@1348_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1349 N_OUT8_Mp8@1349_d N_OUT7_Mp8@1349_g N_VDD_Mp8@1349_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1348 N_OUT8_Mp8@1348_d N_OUT7_Mp8@1348_g N_VDD_Mp8@1348_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1347 N_OUT8_Mn8@1347_d N_OUT7_Mn8@1347_g N_VSS_Mn8@1347_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1346 N_OUT8_Mn8@1346_d N_OUT7_Mn8@1346_g N_VSS_Mn8@1346_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1347 N_OUT8_Mp8@1347_d N_OUT7_Mp8@1347_g N_VDD_Mp8@1347_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1346 N_OUT8_Mp8@1346_d N_OUT7_Mp8@1346_g N_VDD_Mp8@1346_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1345 N_OUT8_Mn8@1345_d N_OUT7_Mn8@1345_g N_VSS_Mn8@1345_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1344 N_OUT8_Mn8@1344_d N_OUT7_Mn8@1344_g N_VSS_Mn8@1344_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1345 N_OUT8_Mp8@1345_d N_OUT7_Mp8@1345_g N_VDD_Mp8@1345_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1344 N_OUT8_Mp8@1344_d N_OUT7_Mp8@1344_g N_VDD_Mp8@1344_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1343 N_OUT8_Mn8@1343_d N_OUT7_Mn8@1343_g N_VSS_Mn8@1343_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1342 N_OUT8_Mn8@1342_d N_OUT7_Mn8@1342_g N_VSS_Mn8@1342_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1343 N_OUT8_Mp8@1343_d N_OUT7_Mp8@1343_g N_VDD_Mp8@1343_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1342 N_OUT8_Mp8@1342_d N_OUT7_Mp8@1342_g N_VDD_Mp8@1342_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1341 N_OUT8_Mn8@1341_d N_OUT7_Mn8@1341_g N_VSS_Mn8@1341_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1340 N_OUT8_Mn8@1340_d N_OUT7_Mn8@1340_g N_VSS_Mn8@1340_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1341 N_OUT8_Mp8@1341_d N_OUT7_Mp8@1341_g N_VDD_Mp8@1341_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1340 N_OUT8_Mp8@1340_d N_OUT7_Mp8@1340_g N_VDD_Mp8@1340_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1339 N_OUT8_Mn8@1339_d N_OUT7_Mn8@1339_g N_VSS_Mn8@1339_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1338 N_OUT8_Mn8@1338_d N_OUT7_Mn8@1338_g N_VSS_Mn8@1338_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1339 N_OUT8_Mp8@1339_d N_OUT7_Mp8@1339_g N_VDD_Mp8@1339_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1338 N_OUT8_Mp8@1338_d N_OUT7_Mp8@1338_g N_VDD_Mp8@1338_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1337 N_OUT8_Mn8@1337_d N_OUT7_Mn8@1337_g N_VSS_Mn8@1337_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1336 N_OUT8_Mn8@1336_d N_OUT7_Mn8@1336_g N_VSS_Mn8@1336_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1337 N_OUT8_Mp8@1337_d N_OUT7_Mp8@1337_g N_VDD_Mp8@1337_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1336 N_OUT8_Mp8@1336_d N_OUT7_Mp8@1336_g N_VDD_Mp8@1336_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1335 N_OUT8_Mn8@1335_d N_OUT7_Mn8@1335_g N_VSS_Mn8@1335_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1334 N_OUT8_Mn8@1334_d N_OUT7_Mn8@1334_g N_VSS_Mn8@1334_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1335 N_OUT8_Mp8@1335_d N_OUT7_Mp8@1335_g N_VDD_Mp8@1335_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1334 N_OUT8_Mp8@1334_d N_OUT7_Mp8@1334_g N_VDD_Mp8@1334_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1333 N_OUT8_Mn8@1333_d N_OUT7_Mn8@1333_g N_VSS_Mn8@1333_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1332 N_OUT8_Mn8@1332_d N_OUT7_Mn8@1332_g N_VSS_Mn8@1332_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1333 N_OUT8_Mp8@1333_d N_OUT7_Mp8@1333_g N_VDD_Mp8@1333_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1332 N_OUT8_Mp8@1332_d N_OUT7_Mp8@1332_g N_VDD_Mp8@1332_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1331 N_OUT8_Mn8@1331_d N_OUT7_Mn8@1331_g N_VSS_Mn8@1331_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1330 N_OUT8_Mn8@1330_d N_OUT7_Mn8@1330_g N_VSS_Mn8@1330_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1331 N_OUT8_Mp8@1331_d N_OUT7_Mp8@1331_g N_VDD_Mp8@1331_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1330 N_OUT8_Mp8@1330_d N_OUT7_Mp8@1330_g N_VDD_Mp8@1330_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1329 N_OUT8_Mn8@1329_d N_OUT7_Mn8@1329_g N_VSS_Mn8@1329_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1328 N_OUT8_Mn8@1328_d N_OUT7_Mn8@1328_g N_VSS_Mn8@1328_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1329 N_OUT8_Mp8@1329_d N_OUT7_Mp8@1329_g N_VDD_Mp8@1329_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1328 N_OUT8_Mp8@1328_d N_OUT7_Mp8@1328_g N_VDD_Mp8@1328_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1327 N_OUT8_Mn8@1327_d N_OUT7_Mn8@1327_g N_VSS_Mn8@1327_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1326 N_OUT8_Mn8@1326_d N_OUT7_Mn8@1326_g N_VSS_Mn8@1326_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1327 N_OUT8_Mp8@1327_d N_OUT7_Mp8@1327_g N_VDD_Mp8@1327_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1326 N_OUT8_Mp8@1326_d N_OUT7_Mp8@1326_g N_VDD_Mp8@1326_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1325 N_OUT8_Mn8@1325_d N_OUT7_Mn8@1325_g N_VSS_Mn8@1325_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1324 N_OUT8_Mn8@1324_d N_OUT7_Mn8@1324_g N_VSS_Mn8@1324_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1325 N_OUT8_Mp8@1325_d N_OUT7_Mp8@1325_g N_VDD_Mp8@1325_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1324 N_OUT8_Mp8@1324_d N_OUT7_Mp8@1324_g N_VDD_Mp8@1324_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1323 N_OUT8_Mn8@1323_d N_OUT7_Mn8@1323_g N_VSS_Mn8@1323_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1322 N_OUT8_Mn8@1322_d N_OUT7_Mn8@1322_g N_VSS_Mn8@1322_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1323 N_OUT8_Mp8@1323_d N_OUT7_Mp8@1323_g N_VDD_Mp8@1323_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1322 N_OUT8_Mp8@1322_d N_OUT7_Mp8@1322_g N_VDD_Mp8@1322_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1321 N_OUT8_Mn8@1321_d N_OUT7_Mn8@1321_g N_VSS_Mn8@1321_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1320 N_OUT8_Mn8@1320_d N_OUT7_Mn8@1320_g N_VSS_Mn8@1320_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1321 N_OUT8_Mp8@1321_d N_OUT7_Mp8@1321_g N_VDD_Mp8@1321_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1320 N_OUT8_Mp8@1320_d N_OUT7_Mp8@1320_g N_VDD_Mp8@1320_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1319 N_OUT8_Mn8@1319_d N_OUT7_Mn8@1319_g N_VSS_Mn8@1319_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1318 N_OUT8_Mn8@1318_d N_OUT7_Mn8@1318_g N_VSS_Mn8@1318_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1319 N_OUT8_Mp8@1319_d N_OUT7_Mp8@1319_g N_VDD_Mp8@1319_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1318 N_OUT8_Mp8@1318_d N_OUT7_Mp8@1318_g N_VDD_Mp8@1318_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1317 N_OUT8_Mn8@1317_d N_OUT7_Mn8@1317_g N_VSS_Mn8@1317_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1316 N_OUT8_Mn8@1316_d N_OUT7_Mn8@1316_g N_VSS_Mn8@1316_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1317 N_OUT8_Mp8@1317_d N_OUT7_Mp8@1317_g N_VDD_Mp8@1317_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1316 N_OUT8_Mp8@1316_d N_OUT7_Mp8@1316_g N_VDD_Mp8@1316_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1315 N_OUT8_Mn8@1315_d N_OUT7_Mn8@1315_g N_VSS_Mn8@1315_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1314 N_OUT8_Mn8@1314_d N_OUT7_Mn8@1314_g N_VSS_Mn8@1314_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1315 N_OUT8_Mp8@1315_d N_OUT7_Mp8@1315_g N_VDD_Mp8@1315_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1314 N_OUT8_Mp8@1314_d N_OUT7_Mp8@1314_g N_VDD_Mp8@1314_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1313 N_OUT8_Mn8@1313_d N_OUT7_Mn8@1313_g N_VSS_Mn8@1313_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1312 N_OUT8_Mn8@1312_d N_OUT7_Mn8@1312_g N_VSS_Mn8@1312_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1313 N_OUT8_Mp8@1313_d N_OUT7_Mp8@1313_g N_VDD_Mp8@1313_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1312 N_OUT8_Mp8@1312_d N_OUT7_Mp8@1312_g N_VDD_Mp8@1312_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1311 N_OUT8_Mn8@1311_d N_OUT7_Mn8@1311_g N_VSS_Mn8@1311_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1310 N_OUT8_Mn8@1310_d N_OUT7_Mn8@1310_g N_VSS_Mn8@1310_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1311 N_OUT8_Mp8@1311_d N_OUT7_Mp8@1311_g N_VDD_Mp8@1311_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1310 N_OUT8_Mp8@1310_d N_OUT7_Mp8@1310_g N_VDD_Mp8@1310_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1309 N_OUT8_Mn8@1309_d N_OUT7_Mn8@1309_g N_VSS_Mn8@1309_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1308 N_OUT8_Mn8@1308_d N_OUT7_Mn8@1308_g N_VSS_Mn8@1308_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1309 N_OUT8_Mp8@1309_d N_OUT7_Mp8@1309_g N_VDD_Mp8@1309_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1308 N_OUT8_Mp8@1308_d N_OUT7_Mp8@1308_g N_VDD_Mp8@1308_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1307 N_OUT8_Mn8@1307_d N_OUT7_Mn8@1307_g N_VSS_Mn8@1307_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1306 N_OUT8_Mn8@1306_d N_OUT7_Mn8@1306_g N_VSS_Mn8@1306_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1307 N_OUT8_Mp8@1307_d N_OUT7_Mp8@1307_g N_VDD_Mp8@1307_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1306 N_OUT8_Mp8@1306_d N_OUT7_Mp8@1306_g N_VDD_Mp8@1306_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1305 N_OUT8_Mn8@1305_d N_OUT7_Mn8@1305_g N_VSS_Mn8@1305_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1304 N_OUT8_Mn8@1304_d N_OUT7_Mn8@1304_g N_VSS_Mn8@1304_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1305 N_OUT8_Mp8@1305_d N_OUT7_Mp8@1305_g N_VDD_Mp8@1305_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1304 N_OUT8_Mp8@1304_d N_OUT7_Mp8@1304_g N_VDD_Mp8@1304_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1303 N_OUT8_Mn8@1303_d N_OUT7_Mn8@1303_g N_VSS_Mn8@1303_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1302 N_OUT8_Mn8@1302_d N_OUT7_Mn8@1302_g N_VSS_Mn8@1302_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1303 N_OUT8_Mp8@1303_d N_OUT7_Mp8@1303_g N_VDD_Mp8@1303_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1302 N_OUT8_Mp8@1302_d N_OUT7_Mp8@1302_g N_VDD_Mp8@1302_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1301 N_OUT8_Mn8@1301_d N_OUT7_Mn8@1301_g N_VSS_Mn8@1301_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1300 N_OUT8_Mn8@1300_d N_OUT7_Mn8@1300_g N_VSS_Mn8@1300_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1301 N_OUT8_Mp8@1301_d N_OUT7_Mp8@1301_g N_VDD_Mp8@1301_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1300 N_OUT8_Mp8@1300_d N_OUT7_Mp8@1300_g N_VDD_Mp8@1300_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1299 N_OUT8_Mn8@1299_d N_OUT7_Mn8@1299_g N_VSS_Mn8@1299_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1298 N_OUT8_Mn8@1298_d N_OUT7_Mn8@1298_g N_VSS_Mn8@1298_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1299 N_OUT8_Mp8@1299_d N_OUT7_Mp8@1299_g N_VDD_Mp8@1299_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1298 N_OUT8_Mp8@1298_d N_OUT7_Mp8@1298_g N_VDD_Mp8@1298_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1297 N_OUT8_Mn8@1297_d N_OUT7_Mn8@1297_g N_VSS_Mn8@1297_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1296 N_OUT8_Mn8@1296_d N_OUT7_Mn8@1296_g N_VSS_Mn8@1296_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1297 N_OUT8_Mp8@1297_d N_OUT7_Mp8@1297_g N_VDD_Mp8@1297_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1296 N_OUT8_Mp8@1296_d N_OUT7_Mp8@1296_g N_VDD_Mp8@1296_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1295 N_OUT8_Mn8@1295_d N_OUT7_Mn8@1295_g N_VSS_Mn8@1295_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1294 N_OUT8_Mn8@1294_d N_OUT7_Mn8@1294_g N_VSS_Mn8@1294_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1295 N_OUT8_Mp8@1295_d N_OUT7_Mp8@1295_g N_VDD_Mp8@1295_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1294 N_OUT8_Mp8@1294_d N_OUT7_Mp8@1294_g N_VDD_Mp8@1294_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1293 N_OUT8_Mn8@1293_d N_OUT7_Mn8@1293_g N_VSS_Mn8@1293_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1292 N_OUT8_Mn8@1292_d N_OUT7_Mn8@1292_g N_VSS_Mn8@1292_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1293 N_OUT8_Mp8@1293_d N_OUT7_Mp8@1293_g N_VDD_Mp8@1293_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1292 N_OUT8_Mp8@1292_d N_OUT7_Mp8@1292_g N_VDD_Mp8@1292_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1291 N_OUT8_Mn8@1291_d N_OUT7_Mn8@1291_g N_VSS_Mn8@1291_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1290 N_OUT8_Mn8@1290_d N_OUT7_Mn8@1290_g N_VSS_Mn8@1290_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1291 N_OUT8_Mp8@1291_d N_OUT7_Mp8@1291_g N_VDD_Mp8@1291_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1290 N_OUT8_Mp8@1290_d N_OUT7_Mp8@1290_g N_VDD_Mp8@1290_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1289 N_OUT8_Mn8@1289_d N_OUT7_Mn8@1289_g N_VSS_Mn8@1289_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1288 N_OUT8_Mn8@1288_d N_OUT7_Mn8@1288_g N_VSS_Mn8@1288_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1289 N_OUT8_Mp8@1289_d N_OUT7_Mp8@1289_g N_VDD_Mp8@1289_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1288 N_OUT8_Mp8@1288_d N_OUT7_Mp8@1288_g N_VDD_Mp8@1288_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1287 N_OUT8_Mn8@1287_d N_OUT7_Mn8@1287_g N_VSS_Mn8@1287_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1286 N_OUT8_Mn8@1286_d N_OUT7_Mn8@1286_g N_VSS_Mn8@1286_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1287 N_OUT8_Mp8@1287_d N_OUT7_Mp8@1287_g N_VDD_Mp8@1287_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1286 N_OUT8_Mp8@1286_d N_OUT7_Mp8@1286_g N_VDD_Mp8@1286_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1285 N_OUT8_Mn8@1285_d N_OUT7_Mn8@1285_g N_VSS_Mn8@1285_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1284 N_OUT8_Mn8@1284_d N_OUT7_Mn8@1284_g N_VSS_Mn8@1284_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1285 N_OUT8_Mp8@1285_d N_OUT7_Mp8@1285_g N_VDD_Mp8@1285_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1284 N_OUT8_Mp8@1284_d N_OUT7_Mp8@1284_g N_VDD_Mp8@1284_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1283 N_OUT8_Mn8@1283_d N_OUT7_Mn8@1283_g N_VSS_Mn8@1283_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1282 N_OUT8_Mn8@1282_d N_OUT7_Mn8@1282_g N_VSS_Mn8@1282_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1283 N_OUT8_Mp8@1283_d N_OUT7_Mp8@1283_g N_VDD_Mp8@1283_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1282 N_OUT8_Mp8@1282_d N_OUT7_Mp8@1282_g N_VDD_Mp8@1282_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1281 N_OUT8_Mn8@1281_d N_OUT7_Mn8@1281_g N_VSS_Mn8@1281_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1280 N_OUT8_Mn8@1280_d N_OUT7_Mn8@1280_g N_VSS_Mn8@1280_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1281 N_OUT8_Mp8@1281_d N_OUT7_Mp8@1281_g N_VDD_Mp8@1281_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1280 N_OUT8_Mp8@1280_d N_OUT7_Mp8@1280_g N_VDD_Mp8@1280_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1279 N_OUT8_Mn8@1279_d N_OUT7_Mn8@1279_g N_VSS_Mn8@1279_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1278 N_OUT8_Mn8@1278_d N_OUT7_Mn8@1278_g N_VSS_Mn8@1278_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1279 N_OUT8_Mp8@1279_d N_OUT7_Mp8@1279_g N_VDD_Mp8@1279_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1278 N_OUT8_Mp8@1278_d N_OUT7_Mp8@1278_g N_VDD_Mp8@1278_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1277 N_OUT8_Mn8@1277_d N_OUT7_Mn8@1277_g N_VSS_Mn8@1277_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1276 N_OUT8_Mn8@1276_d N_OUT7_Mn8@1276_g N_VSS_Mn8@1276_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1277 N_OUT8_Mp8@1277_d N_OUT7_Mp8@1277_g N_VDD_Mp8@1277_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1276 N_OUT8_Mp8@1276_d N_OUT7_Mp8@1276_g N_VDD_Mp8@1276_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1275 N_OUT8_Mn8@1275_d N_OUT7_Mn8@1275_g N_VSS_Mn8@1275_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1274 N_OUT8_Mn8@1274_d N_OUT7_Mn8@1274_g N_VSS_Mn8@1274_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1275 N_OUT8_Mp8@1275_d N_OUT7_Mp8@1275_g N_VDD_Mp8@1275_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1274 N_OUT8_Mp8@1274_d N_OUT7_Mp8@1274_g N_VDD_Mp8@1274_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1273 N_OUT8_Mn8@1273_d N_OUT7_Mn8@1273_g N_VSS_Mn8@1273_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1272 N_OUT8_Mn8@1272_d N_OUT7_Mn8@1272_g N_VSS_Mn8@1272_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1273 N_OUT8_Mp8@1273_d N_OUT7_Mp8@1273_g N_VDD_Mp8@1273_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1272 N_OUT8_Mp8@1272_d N_OUT7_Mp8@1272_g N_VDD_Mp8@1272_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1271 N_OUT8_Mn8@1271_d N_OUT7_Mn8@1271_g N_VSS_Mn8@1271_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1270 N_OUT8_Mn8@1270_d N_OUT7_Mn8@1270_g N_VSS_Mn8@1270_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1271 N_OUT8_Mp8@1271_d N_OUT7_Mp8@1271_g N_VDD_Mp8@1271_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1270 N_OUT8_Mp8@1270_d N_OUT7_Mp8@1270_g N_VDD_Mp8@1270_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1269 N_OUT8_Mn8@1269_d N_OUT7_Mn8@1269_g N_VSS_Mn8@1269_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1268 N_OUT8_Mn8@1268_d N_OUT7_Mn8@1268_g N_VSS_Mn8@1268_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1269 N_OUT8_Mp8@1269_d N_OUT7_Mp8@1269_g N_VDD_Mp8@1269_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1268 N_OUT8_Mp8@1268_d N_OUT7_Mp8@1268_g N_VDD_Mp8@1268_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1267 N_OUT8_Mn8@1267_d N_OUT7_Mn8@1267_g N_VSS_Mn8@1267_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1266 N_OUT8_Mn8@1266_d N_OUT7_Mn8@1266_g N_VSS_Mn8@1266_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1267 N_OUT8_Mp8@1267_d N_OUT7_Mp8@1267_g N_VDD_Mp8@1267_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1266 N_OUT8_Mp8@1266_d N_OUT7_Mp8@1266_g N_VDD_Mp8@1266_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1265 N_OUT8_Mn8@1265_d N_OUT7_Mn8@1265_g N_VSS_Mn8@1265_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1264 N_OUT8_Mn8@1264_d N_OUT7_Mn8@1264_g N_VSS_Mn8@1264_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1265 N_OUT8_Mp8@1265_d N_OUT7_Mp8@1265_g N_VDD_Mp8@1265_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1264 N_OUT8_Mp8@1264_d N_OUT7_Mp8@1264_g N_VDD_Mp8@1264_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1263 N_OUT8_Mn8@1263_d N_OUT7_Mn8@1263_g N_VSS_Mn8@1263_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1262 N_OUT8_Mn8@1262_d N_OUT7_Mn8@1262_g N_VSS_Mn8@1262_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1263 N_OUT8_Mp8@1263_d N_OUT7_Mp8@1263_g N_VDD_Mp8@1263_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1262 N_OUT8_Mp8@1262_d N_OUT7_Mp8@1262_g N_VDD_Mp8@1262_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1261 N_OUT8_Mn8@1261_d N_OUT7_Mn8@1261_g N_VSS_Mn8@1261_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1260 N_OUT8_Mn8@1260_d N_OUT7_Mn8@1260_g N_VSS_Mn8@1260_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1261 N_OUT8_Mp8@1261_d N_OUT7_Mp8@1261_g N_VDD_Mp8@1261_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1260 N_OUT8_Mp8@1260_d N_OUT7_Mp8@1260_g N_VDD_Mp8@1260_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1259 N_OUT8_Mn8@1259_d N_OUT7_Mn8@1259_g N_VSS_Mn8@1259_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1258 N_OUT8_Mn8@1258_d N_OUT7_Mn8@1258_g N_VSS_Mn8@1258_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1259 N_OUT8_Mp8@1259_d N_OUT7_Mp8@1259_g N_VDD_Mp8@1259_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1258 N_OUT8_Mp8@1258_d N_OUT7_Mp8@1258_g N_VDD_Mp8@1258_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1257 N_OUT8_Mn8@1257_d N_OUT7_Mn8@1257_g N_VSS_Mn8@1257_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1256 N_OUT8_Mn8@1256_d N_OUT7_Mn8@1256_g N_VSS_Mn8@1256_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1257 N_OUT8_Mp8@1257_d N_OUT7_Mp8@1257_g N_VDD_Mp8@1257_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1256 N_OUT8_Mp8@1256_d N_OUT7_Mp8@1256_g N_VDD_Mp8@1256_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1255 N_OUT8_Mn8@1255_d N_OUT7_Mn8@1255_g N_VSS_Mn8@1255_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1254 N_OUT8_Mn8@1254_d N_OUT7_Mn8@1254_g N_VSS_Mn8@1254_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1255 N_OUT8_Mp8@1255_d N_OUT7_Mp8@1255_g N_VDD_Mp8@1255_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1254 N_OUT8_Mp8@1254_d N_OUT7_Mp8@1254_g N_VDD_Mp8@1254_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1253 N_OUT8_Mn8@1253_d N_OUT7_Mn8@1253_g N_VSS_Mn8@1253_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1252 N_OUT8_Mn8@1252_d N_OUT7_Mn8@1252_g N_VSS_Mn8@1252_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1253 N_OUT8_Mp8@1253_d N_OUT7_Mp8@1253_g N_VDD_Mp8@1253_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1252 N_OUT8_Mp8@1252_d N_OUT7_Mp8@1252_g N_VDD_Mp8@1252_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1251 N_OUT8_Mn8@1251_d N_OUT7_Mn8@1251_g N_VSS_Mn8@1251_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1250 N_OUT8_Mn8@1250_d N_OUT7_Mn8@1250_g N_VSS_Mn8@1250_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1251 N_OUT8_Mp8@1251_d N_OUT7_Mp8@1251_g N_VDD_Mp8@1251_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1250 N_OUT8_Mp8@1250_d N_OUT7_Mp8@1250_g N_VDD_Mp8@1250_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1249 N_OUT8_Mn8@1249_d N_OUT7_Mn8@1249_g N_VSS_Mn8@1249_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1248 N_OUT8_Mn8@1248_d N_OUT7_Mn8@1248_g N_VSS_Mn8@1248_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1249 N_OUT8_Mp8@1249_d N_OUT7_Mp8@1249_g N_VDD_Mp8@1249_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1248 N_OUT8_Mp8@1248_d N_OUT7_Mp8@1248_g N_VDD_Mp8@1248_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1247 N_OUT8_Mn8@1247_d N_OUT7_Mn8@1247_g N_VSS_Mn8@1247_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1246 N_OUT8_Mn8@1246_d N_OUT7_Mn8@1246_g N_VSS_Mn8@1246_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1247 N_OUT8_Mp8@1247_d N_OUT7_Mp8@1247_g N_VDD_Mp8@1247_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1246 N_OUT8_Mp8@1246_d N_OUT7_Mp8@1246_g N_VDD_Mp8@1246_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1245 N_OUT8_Mn8@1245_d N_OUT7_Mn8@1245_g N_VSS_Mn8@1245_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1244 N_OUT8_Mn8@1244_d N_OUT7_Mn8@1244_g N_VSS_Mn8@1244_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1245 N_OUT8_Mp8@1245_d N_OUT7_Mp8@1245_g N_VDD_Mp8@1245_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1244 N_OUT8_Mp8@1244_d N_OUT7_Mp8@1244_g N_VDD_Mp8@1244_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1243 N_OUT8_Mn8@1243_d N_OUT7_Mn8@1243_g N_VSS_Mn8@1243_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1242 N_OUT8_Mn8@1242_d N_OUT7_Mn8@1242_g N_VSS_Mn8@1242_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1243 N_OUT8_Mp8@1243_d N_OUT7_Mp8@1243_g N_VDD_Mp8@1243_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1242 N_OUT8_Mp8@1242_d N_OUT7_Mp8@1242_g N_VDD_Mp8@1242_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1241 N_OUT8_Mn8@1241_d N_OUT7_Mn8@1241_g N_VSS_Mn8@1241_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1240 N_OUT8_Mn8@1240_d N_OUT7_Mn8@1240_g N_VSS_Mn8@1240_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1241 N_OUT8_Mp8@1241_d N_OUT7_Mp8@1241_g N_VDD_Mp8@1241_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1240 N_OUT8_Mp8@1240_d N_OUT7_Mp8@1240_g N_VDD_Mp8@1240_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1239 N_OUT8_Mn8@1239_d N_OUT7_Mn8@1239_g N_VSS_Mn8@1239_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1238 N_OUT8_Mn8@1238_d N_OUT7_Mn8@1238_g N_VSS_Mn8@1238_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1239 N_OUT8_Mp8@1239_d N_OUT7_Mp8@1239_g N_VDD_Mp8@1239_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1238 N_OUT8_Mp8@1238_d N_OUT7_Mp8@1238_g N_VDD_Mp8@1238_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1237 N_OUT8_Mn8@1237_d N_OUT7_Mn8@1237_g N_VSS_Mn8@1237_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1236 N_OUT8_Mn8@1236_d N_OUT7_Mn8@1236_g N_VSS_Mn8@1236_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1237 N_OUT8_Mp8@1237_d N_OUT7_Mp8@1237_g N_VDD_Mp8@1237_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1236 N_OUT8_Mp8@1236_d N_OUT7_Mp8@1236_g N_VDD_Mp8@1236_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1235 N_OUT8_Mn8@1235_d N_OUT7_Mn8@1235_g N_VSS_Mn8@1235_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1234 N_OUT8_Mn8@1234_d N_OUT7_Mn8@1234_g N_VSS_Mn8@1234_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1235 N_OUT8_Mp8@1235_d N_OUT7_Mp8@1235_g N_VDD_Mp8@1235_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1234 N_OUT8_Mp8@1234_d N_OUT7_Mp8@1234_g N_VDD_Mp8@1234_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1233 N_OUT8_Mn8@1233_d N_OUT7_Mn8@1233_g N_VSS_Mn8@1233_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1232 N_OUT8_Mn8@1232_d N_OUT7_Mn8@1232_g N_VSS_Mn8@1232_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1233 N_OUT8_Mp8@1233_d N_OUT7_Mp8@1233_g N_VDD_Mp8@1233_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1232 N_OUT8_Mp8@1232_d N_OUT7_Mp8@1232_g N_VDD_Mp8@1232_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1231 N_OUT8_Mn8@1231_d N_OUT7_Mn8@1231_g N_VSS_Mn8@1231_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1230 N_OUT8_Mn8@1230_d N_OUT7_Mn8@1230_g N_VSS_Mn8@1230_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1231 N_OUT8_Mp8@1231_d N_OUT7_Mp8@1231_g N_VDD_Mp8@1231_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1230 N_OUT8_Mp8@1230_d N_OUT7_Mp8@1230_g N_VDD_Mp8@1230_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1229 N_OUT8_Mn8@1229_d N_OUT7_Mn8@1229_g N_VSS_Mn8@1229_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1228 N_OUT8_Mn8@1228_d N_OUT7_Mn8@1228_g N_VSS_Mn8@1228_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1229 N_OUT8_Mp8@1229_d N_OUT7_Mp8@1229_g N_VDD_Mp8@1229_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1228 N_OUT8_Mp8@1228_d N_OUT7_Mp8@1228_g N_VDD_Mp8@1228_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1227 N_OUT8_Mn8@1227_d N_OUT7_Mn8@1227_g N_VSS_Mn8@1227_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1226 N_OUT8_Mn8@1226_d N_OUT7_Mn8@1226_g N_VSS_Mn8@1226_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1227 N_OUT8_Mp8@1227_d N_OUT7_Mp8@1227_g N_VDD_Mp8@1227_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1226 N_OUT8_Mp8@1226_d N_OUT7_Mp8@1226_g N_VDD_Mp8@1226_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1225 N_OUT8_Mn8@1225_d N_OUT7_Mn8@1225_g N_VSS_Mn8@1225_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1224 N_OUT8_Mn8@1224_d N_OUT7_Mn8@1224_g N_VSS_Mn8@1224_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1225 N_OUT8_Mp8@1225_d N_OUT7_Mp8@1225_g N_VDD_Mp8@1225_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1224 N_OUT8_Mp8@1224_d N_OUT7_Mp8@1224_g N_VDD_Mp8@1224_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1223 N_OUT8_Mn8@1223_d N_OUT7_Mn8@1223_g N_VSS_Mn8@1223_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1222 N_OUT8_Mn8@1222_d N_OUT7_Mn8@1222_g N_VSS_Mn8@1222_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1223 N_OUT8_Mp8@1223_d N_OUT7_Mp8@1223_g N_VDD_Mp8@1223_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1222 N_OUT8_Mp8@1222_d N_OUT7_Mp8@1222_g N_VDD_Mp8@1222_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1221 N_OUT8_Mn8@1221_d N_OUT7_Mn8@1221_g N_VSS_Mn8@1221_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1220 N_OUT8_Mn8@1220_d N_OUT7_Mn8@1220_g N_VSS_Mn8@1220_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1221 N_OUT8_Mp8@1221_d N_OUT7_Mp8@1221_g N_VDD_Mp8@1221_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1220 N_OUT8_Mp8@1220_d N_OUT7_Mp8@1220_g N_VDD_Mp8@1220_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1219 N_OUT8_Mn8@1219_d N_OUT7_Mn8@1219_g N_VSS_Mn8@1219_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1218 N_OUT8_Mn8@1218_d N_OUT7_Mn8@1218_g N_VSS_Mn8@1218_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1219 N_OUT8_Mp8@1219_d N_OUT7_Mp8@1219_g N_VDD_Mp8@1219_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1218 N_OUT8_Mp8@1218_d N_OUT7_Mp8@1218_g N_VDD_Mp8@1218_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1217 N_OUT8_Mn8@1217_d N_OUT7_Mn8@1217_g N_VSS_Mn8@1217_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1216 N_OUT8_Mn8@1216_d N_OUT7_Mn8@1216_g N_VSS_Mn8@1216_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1217 N_OUT8_Mp8@1217_d N_OUT7_Mp8@1217_g N_VDD_Mp8@1217_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1216 N_OUT8_Mp8@1216_d N_OUT7_Mp8@1216_g N_VDD_Mp8@1216_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1215 N_OUT8_Mn8@1215_d N_OUT7_Mn8@1215_g N_VSS_Mn8@1215_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1214 N_OUT8_Mn8@1214_d N_OUT7_Mn8@1214_g N_VSS_Mn8@1214_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1215 N_OUT8_Mp8@1215_d N_OUT7_Mp8@1215_g N_VDD_Mp8@1215_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1214 N_OUT8_Mp8@1214_d N_OUT7_Mp8@1214_g N_VDD_Mp8@1214_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1213 N_OUT8_Mn8@1213_d N_OUT7_Mn8@1213_g N_VSS_Mn8@1213_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1212 N_OUT8_Mn8@1212_d N_OUT7_Mn8@1212_g N_VSS_Mn8@1212_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1213 N_OUT8_Mp8@1213_d N_OUT7_Mp8@1213_g N_VDD_Mp8@1213_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1212 N_OUT8_Mp8@1212_d N_OUT7_Mp8@1212_g N_VDD_Mp8@1212_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1211 N_OUT8_Mn8@1211_d N_OUT7_Mn8@1211_g N_VSS_Mn8@1211_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1210 N_OUT8_Mn8@1210_d N_OUT7_Mn8@1210_g N_VSS_Mn8@1210_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1211 N_OUT8_Mp8@1211_d N_OUT7_Mp8@1211_g N_VDD_Mp8@1211_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1210 N_OUT8_Mp8@1210_d N_OUT7_Mp8@1210_g N_VDD_Mp8@1210_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1209 N_OUT8_Mn8@1209_d N_OUT7_Mn8@1209_g N_VSS_Mn8@1209_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1208 N_OUT8_Mn8@1208_d N_OUT7_Mn8@1208_g N_VSS_Mn8@1208_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1209 N_OUT8_Mp8@1209_d N_OUT7_Mp8@1209_g N_VDD_Mp8@1209_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1208 N_OUT8_Mp8@1208_d N_OUT7_Mp8@1208_g N_VDD_Mp8@1208_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1207 N_OUT8_Mn8@1207_d N_OUT7_Mn8@1207_g N_VSS_Mn8@1207_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1206 N_OUT8_Mn8@1206_d N_OUT7_Mn8@1206_g N_VSS_Mn8@1206_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1207 N_OUT8_Mp8@1207_d N_OUT7_Mp8@1207_g N_VDD_Mp8@1207_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1206 N_OUT8_Mp8@1206_d N_OUT7_Mp8@1206_g N_VDD_Mp8@1206_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1205 N_OUT8_Mn8@1205_d N_OUT7_Mn8@1205_g N_VSS_Mn8@1205_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1204 N_OUT8_Mn8@1204_d N_OUT7_Mn8@1204_g N_VSS_Mn8@1204_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1205 N_OUT8_Mp8@1205_d N_OUT7_Mp8@1205_g N_VDD_Mp8@1205_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1204 N_OUT8_Mp8@1204_d N_OUT7_Mp8@1204_g N_VDD_Mp8@1204_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1203 N_OUT8_Mn8@1203_d N_OUT7_Mn8@1203_g N_VSS_Mn8@1203_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1202 N_OUT8_Mn8@1202_d N_OUT7_Mn8@1202_g N_VSS_Mn8@1202_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1203 N_OUT8_Mp8@1203_d N_OUT7_Mp8@1203_g N_VDD_Mp8@1203_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1202 N_OUT8_Mp8@1202_d N_OUT7_Mp8@1202_g N_VDD_Mp8@1202_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1201 N_OUT8_Mn8@1201_d N_OUT7_Mn8@1201_g N_VSS_Mn8@1201_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1200 N_OUT8_Mn8@1200_d N_OUT7_Mn8@1200_g N_VSS_Mn8@1200_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1201 N_OUT8_Mp8@1201_d N_OUT7_Mp8@1201_g N_VDD_Mp8@1201_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1200 N_OUT8_Mp8@1200_d N_OUT7_Mp8@1200_g N_VDD_Mp8@1200_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1199 N_OUT8_Mn8@1199_d N_OUT7_Mn8@1199_g N_VSS_Mn8@1199_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1198 N_OUT8_Mn8@1198_d N_OUT7_Mn8@1198_g N_VSS_Mn8@1198_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1199 N_OUT8_Mp8@1199_d N_OUT7_Mp8@1199_g N_VDD_Mp8@1199_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1198 N_OUT8_Mp8@1198_d N_OUT7_Mp8@1198_g N_VDD_Mp8@1198_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1197 N_OUT8_Mn8@1197_d N_OUT7_Mn8@1197_g N_VSS_Mn8@1197_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1196 N_OUT8_Mn8@1196_d N_OUT7_Mn8@1196_g N_VSS_Mn8@1196_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1197 N_OUT8_Mp8@1197_d N_OUT7_Mp8@1197_g N_VDD_Mp8@1197_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1196 N_OUT8_Mp8@1196_d N_OUT7_Mp8@1196_g N_VDD_Mp8@1196_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1195 N_OUT8_Mn8@1195_d N_OUT7_Mn8@1195_g N_VSS_Mn8@1195_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1194 N_OUT8_Mn8@1194_d N_OUT7_Mn8@1194_g N_VSS_Mn8@1194_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1195 N_OUT8_Mp8@1195_d N_OUT7_Mp8@1195_g N_VDD_Mp8@1195_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1194 N_OUT8_Mp8@1194_d N_OUT7_Mp8@1194_g N_VDD_Mp8@1194_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1193 N_OUT8_Mn8@1193_d N_OUT7_Mn8@1193_g N_VSS_Mn8@1193_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1192 N_OUT8_Mn8@1192_d N_OUT7_Mn8@1192_g N_VSS_Mn8@1192_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1193 N_OUT8_Mp8@1193_d N_OUT7_Mp8@1193_g N_VDD_Mp8@1193_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1192 N_OUT8_Mp8@1192_d N_OUT7_Mp8@1192_g N_VDD_Mp8@1192_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1191 N_OUT8_Mn8@1191_d N_OUT7_Mn8@1191_g N_VSS_Mn8@1191_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1190 N_OUT8_Mn8@1190_d N_OUT7_Mn8@1190_g N_VSS_Mn8@1190_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1191 N_OUT8_Mp8@1191_d N_OUT7_Mp8@1191_g N_VDD_Mp8@1191_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1190 N_OUT8_Mp8@1190_d N_OUT7_Mp8@1190_g N_VDD_Mp8@1190_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1189 N_OUT8_Mn8@1189_d N_OUT7_Mn8@1189_g N_VSS_Mn8@1189_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1188 N_OUT8_Mn8@1188_d N_OUT7_Mn8@1188_g N_VSS_Mn8@1188_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1189 N_OUT8_Mp8@1189_d N_OUT7_Mp8@1189_g N_VDD_Mp8@1189_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1188 N_OUT8_Mp8@1188_d N_OUT7_Mp8@1188_g N_VDD_Mp8@1188_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1187 N_OUT8_Mn8@1187_d N_OUT7_Mn8@1187_g N_VSS_Mn8@1187_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1186 N_OUT8_Mn8@1186_d N_OUT7_Mn8@1186_g N_VSS_Mn8@1186_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1187 N_OUT8_Mp8@1187_d N_OUT7_Mp8@1187_g N_VDD_Mp8@1187_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1186 N_OUT8_Mp8@1186_d N_OUT7_Mp8@1186_g N_VDD_Mp8@1186_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1185 N_OUT8_Mn8@1185_d N_OUT7_Mn8@1185_g N_VSS_Mn8@1185_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1184 N_OUT8_Mn8@1184_d N_OUT7_Mn8@1184_g N_VSS_Mn8@1184_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1185 N_OUT8_Mp8@1185_d N_OUT7_Mp8@1185_g N_VDD_Mp8@1185_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1184 N_OUT8_Mp8@1184_d N_OUT7_Mp8@1184_g N_VDD_Mp8@1184_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1183 N_OUT8_Mn8@1183_d N_OUT7_Mn8@1183_g N_VSS_Mn8@1183_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1182 N_OUT8_Mn8@1182_d N_OUT7_Mn8@1182_g N_VSS_Mn8@1182_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1183 N_OUT8_Mp8@1183_d N_OUT7_Mp8@1183_g N_VDD_Mp8@1183_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1182 N_OUT8_Mp8@1182_d N_OUT7_Mp8@1182_g N_VDD_Mp8@1182_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1181 N_OUT8_Mn8@1181_d N_OUT7_Mn8@1181_g N_VSS_Mn8@1181_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1180 N_OUT8_Mn8@1180_d N_OUT7_Mn8@1180_g N_VSS_Mn8@1180_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1181 N_OUT8_Mp8@1181_d N_OUT7_Mp8@1181_g N_VDD_Mp8@1181_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1180 N_OUT8_Mp8@1180_d N_OUT7_Mp8@1180_g N_VDD_Mp8@1180_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1179 N_OUT8_Mn8@1179_d N_OUT7_Mn8@1179_g N_VSS_Mn8@1179_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1178 N_OUT8_Mn8@1178_d N_OUT7_Mn8@1178_g N_VSS_Mn8@1178_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1179 N_OUT8_Mp8@1179_d N_OUT7_Mp8@1179_g N_VDD_Mp8@1179_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1178 N_OUT8_Mp8@1178_d N_OUT7_Mp8@1178_g N_VDD_Mp8@1178_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1177 N_OUT8_Mn8@1177_d N_OUT7_Mn8@1177_g N_VSS_Mn8@1177_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1176 N_OUT8_Mn8@1176_d N_OUT7_Mn8@1176_g N_VSS_Mn8@1176_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1177 N_OUT8_Mp8@1177_d N_OUT7_Mp8@1177_g N_VDD_Mp8@1177_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1176 N_OUT8_Mp8@1176_d N_OUT7_Mp8@1176_g N_VDD_Mp8@1176_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1175 N_OUT8_Mn8@1175_d N_OUT7_Mn8@1175_g N_VSS_Mn8@1175_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1174 N_OUT8_Mn8@1174_d N_OUT7_Mn8@1174_g N_VSS_Mn8@1174_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1175 N_OUT8_Mp8@1175_d N_OUT7_Mp8@1175_g N_VDD_Mp8@1175_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1174 N_OUT8_Mp8@1174_d N_OUT7_Mp8@1174_g N_VDD_Mp8@1174_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1173 N_OUT8_Mn8@1173_d N_OUT7_Mn8@1173_g N_VSS_Mn8@1173_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1172 N_OUT8_Mn8@1172_d N_OUT7_Mn8@1172_g N_VSS_Mn8@1172_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1173 N_OUT8_Mp8@1173_d N_OUT7_Mp8@1173_g N_VDD_Mp8@1173_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1172 N_OUT8_Mp8@1172_d N_OUT7_Mp8@1172_g N_VDD_Mp8@1172_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1171 N_OUT8_Mn8@1171_d N_OUT7_Mn8@1171_g N_VSS_Mn8@1171_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1170 N_OUT8_Mn8@1170_d N_OUT7_Mn8@1170_g N_VSS_Mn8@1170_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1171 N_OUT8_Mp8@1171_d N_OUT7_Mp8@1171_g N_VDD_Mp8@1171_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1170 N_OUT8_Mp8@1170_d N_OUT7_Mp8@1170_g N_VDD_Mp8@1170_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1169 N_OUT8_Mn8@1169_d N_OUT7_Mn8@1169_g N_VSS_Mn8@1169_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1168 N_OUT8_Mn8@1168_d N_OUT7_Mn8@1168_g N_VSS_Mn8@1168_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1169 N_OUT8_Mp8@1169_d N_OUT7_Mp8@1169_g N_VDD_Mp8@1169_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1168 N_OUT8_Mp8@1168_d N_OUT7_Mp8@1168_g N_VDD_Mp8@1168_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1167 N_OUT8_Mn8@1167_d N_OUT7_Mn8@1167_g N_VSS_Mn8@1167_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1166 N_OUT8_Mn8@1166_d N_OUT7_Mn8@1166_g N_VSS_Mn8@1166_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1167 N_OUT8_Mp8@1167_d N_OUT7_Mp8@1167_g N_VDD_Mp8@1167_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1166 N_OUT8_Mp8@1166_d N_OUT7_Mp8@1166_g N_VDD_Mp8@1166_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1165 N_OUT8_Mn8@1165_d N_OUT7_Mn8@1165_g N_VSS_Mn8@1165_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1164 N_OUT8_Mn8@1164_d N_OUT7_Mn8@1164_g N_VSS_Mn8@1164_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1165 N_OUT8_Mp8@1165_d N_OUT7_Mp8@1165_g N_VDD_Mp8@1165_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1164 N_OUT8_Mp8@1164_d N_OUT7_Mp8@1164_g N_VDD_Mp8@1164_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1163 N_OUT8_Mn8@1163_d N_OUT7_Mn8@1163_g N_VSS_Mn8@1163_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1162 N_OUT8_Mn8@1162_d N_OUT7_Mn8@1162_g N_VSS_Mn8@1162_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1163 N_OUT8_Mp8@1163_d N_OUT7_Mp8@1163_g N_VDD_Mp8@1163_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1162 N_OUT8_Mp8@1162_d N_OUT7_Mp8@1162_g N_VDD_Mp8@1162_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1161 N_OUT8_Mn8@1161_d N_OUT7_Mn8@1161_g N_VSS_Mn8@1161_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1160 N_OUT8_Mn8@1160_d N_OUT7_Mn8@1160_g N_VSS_Mn8@1160_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1161 N_OUT8_Mp8@1161_d N_OUT7_Mp8@1161_g N_VDD_Mp8@1161_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1160 N_OUT8_Mp8@1160_d N_OUT7_Mp8@1160_g N_VDD_Mp8@1160_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1159 N_OUT8_Mn8@1159_d N_OUT7_Mn8@1159_g N_VSS_Mn8@1159_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1158 N_OUT8_Mn8@1158_d N_OUT7_Mn8@1158_g N_VSS_Mn8@1158_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1159 N_OUT8_Mp8@1159_d N_OUT7_Mp8@1159_g N_VDD_Mp8@1159_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1158 N_OUT8_Mp8@1158_d N_OUT7_Mp8@1158_g N_VDD_Mp8@1158_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1157 N_OUT8_Mn8@1157_d N_OUT7_Mn8@1157_g N_VSS_Mn8@1157_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1156 N_OUT8_Mn8@1156_d N_OUT7_Mn8@1156_g N_VSS_Mn8@1156_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1157 N_OUT8_Mp8@1157_d N_OUT7_Mp8@1157_g N_VDD_Mp8@1157_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1156 N_OUT8_Mp8@1156_d N_OUT7_Mp8@1156_g N_VDD_Mp8@1156_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1155 N_OUT8_Mn8@1155_d N_OUT7_Mn8@1155_g N_VSS_Mn8@1155_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1154 N_OUT8_Mn8@1154_d N_OUT7_Mn8@1154_g N_VSS_Mn8@1154_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1155 N_OUT8_Mp8@1155_d N_OUT7_Mp8@1155_g N_VDD_Mp8@1155_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1154 N_OUT8_Mp8@1154_d N_OUT7_Mp8@1154_g N_VDD_Mp8@1154_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1153 N_OUT8_Mn8@1153_d N_OUT7_Mn8@1153_g N_VSS_Mn8@1153_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1152 N_OUT8_Mn8@1152_d N_OUT7_Mn8@1152_g N_VSS_Mn8@1152_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1153 N_OUT8_Mp8@1153_d N_OUT7_Mp8@1153_g N_VDD_Mp8@1153_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1152 N_OUT8_Mp8@1152_d N_OUT7_Mp8@1152_g N_VDD_Mp8@1152_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1151 N_OUT8_Mn8@1151_d N_OUT7_Mn8@1151_g N_VSS_Mn8@1151_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1150 N_OUT8_Mn8@1150_d N_OUT7_Mn8@1150_g N_VSS_Mn8@1150_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1151 N_OUT8_Mp8@1151_d N_OUT7_Mp8@1151_g N_VDD_Mp8@1151_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1150 N_OUT8_Mp8@1150_d N_OUT7_Mp8@1150_g N_VDD_Mp8@1150_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1149 N_OUT8_Mn8@1149_d N_OUT7_Mn8@1149_g N_VSS_Mn8@1149_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1148 N_OUT8_Mn8@1148_d N_OUT7_Mn8@1148_g N_VSS_Mn8@1148_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1149 N_OUT8_Mp8@1149_d N_OUT7_Mp8@1149_g N_VDD_Mp8@1149_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1148 N_OUT8_Mp8@1148_d N_OUT7_Mp8@1148_g N_VDD_Mp8@1148_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1147 N_OUT8_Mn8@1147_d N_OUT7_Mn8@1147_g N_VSS_Mn8@1147_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1146 N_OUT8_Mn8@1146_d N_OUT7_Mn8@1146_g N_VSS_Mn8@1146_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1147 N_OUT8_Mp8@1147_d N_OUT7_Mp8@1147_g N_VDD_Mp8@1147_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1146 N_OUT8_Mp8@1146_d N_OUT7_Mp8@1146_g N_VDD_Mp8@1146_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1145 N_OUT8_Mn8@1145_d N_OUT7_Mn8@1145_g N_VSS_Mn8@1145_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1144 N_OUT8_Mn8@1144_d N_OUT7_Mn8@1144_g N_VSS_Mn8@1144_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1145 N_OUT8_Mp8@1145_d N_OUT7_Mp8@1145_g N_VDD_Mp8@1145_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1144 N_OUT8_Mp8@1144_d N_OUT7_Mp8@1144_g N_VDD_Mp8@1144_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1143 N_OUT8_Mn8@1143_d N_OUT7_Mn8@1143_g N_VSS_Mn8@1143_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1142 N_OUT8_Mn8@1142_d N_OUT7_Mn8@1142_g N_VSS_Mn8@1142_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1143 N_OUT8_Mp8@1143_d N_OUT7_Mp8@1143_g N_VDD_Mp8@1143_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1142 N_OUT8_Mp8@1142_d N_OUT7_Mp8@1142_g N_VDD_Mp8@1142_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1141 N_OUT8_Mn8@1141_d N_OUT7_Mn8@1141_g N_VSS_Mn8@1141_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1140 N_OUT8_Mn8@1140_d N_OUT7_Mn8@1140_g N_VSS_Mn8@1140_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1141 N_OUT8_Mp8@1141_d N_OUT7_Mp8@1141_g N_VDD_Mp8@1141_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1140 N_OUT8_Mp8@1140_d N_OUT7_Mp8@1140_g N_VDD_Mp8@1140_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1139 N_OUT8_Mn8@1139_d N_OUT7_Mn8@1139_g N_VSS_Mn8@1139_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1138 N_OUT8_Mn8@1138_d N_OUT7_Mn8@1138_g N_VSS_Mn8@1138_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1139 N_OUT8_Mp8@1139_d N_OUT7_Mp8@1139_g N_VDD_Mp8@1139_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1138 N_OUT8_Mp8@1138_d N_OUT7_Mp8@1138_g N_VDD_Mp8@1138_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1137 N_OUT8_Mn8@1137_d N_OUT7_Mn8@1137_g N_VSS_Mn8@1137_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1136 N_OUT8_Mn8@1136_d N_OUT7_Mn8@1136_g N_VSS_Mn8@1136_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1137 N_OUT8_Mp8@1137_d N_OUT7_Mp8@1137_g N_VDD_Mp8@1137_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1136 N_OUT8_Mp8@1136_d N_OUT7_Mp8@1136_g N_VDD_Mp8@1136_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1135 N_OUT8_Mn8@1135_d N_OUT7_Mn8@1135_g N_VSS_Mn8@1135_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1134 N_OUT8_Mn8@1134_d N_OUT7_Mn8@1134_g N_VSS_Mn8@1134_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1135 N_OUT8_Mp8@1135_d N_OUT7_Mp8@1135_g N_VDD_Mp8@1135_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1134 N_OUT8_Mp8@1134_d N_OUT7_Mp8@1134_g N_VDD_Mp8@1134_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1133 N_OUT8_Mn8@1133_d N_OUT7_Mn8@1133_g N_VSS_Mn8@1133_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1132 N_OUT8_Mn8@1132_d N_OUT7_Mn8@1132_g N_VSS_Mn8@1132_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1133 N_OUT8_Mp8@1133_d N_OUT7_Mp8@1133_g N_VDD_Mp8@1133_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1132 N_OUT8_Mp8@1132_d N_OUT7_Mp8@1132_g N_VDD_Mp8@1132_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1131 N_OUT8_Mn8@1131_d N_OUT7_Mn8@1131_g N_VSS_Mn8@1131_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1130 N_OUT8_Mn8@1130_d N_OUT7_Mn8@1130_g N_VSS_Mn8@1130_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1131 N_OUT8_Mp8@1131_d N_OUT7_Mp8@1131_g N_VDD_Mp8@1131_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1130 N_OUT8_Mp8@1130_d N_OUT7_Mp8@1130_g N_VDD_Mp8@1130_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1129 N_OUT8_Mn8@1129_d N_OUT7_Mn8@1129_g N_VSS_Mn8@1129_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1128 N_OUT8_Mn8@1128_d N_OUT7_Mn8@1128_g N_VSS_Mn8@1128_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1129 N_OUT8_Mp8@1129_d N_OUT7_Mp8@1129_g N_VDD_Mp8@1129_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1128 N_OUT8_Mp8@1128_d N_OUT7_Mp8@1128_g N_VDD_Mp8@1128_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1127 N_OUT8_Mn8@1127_d N_OUT7_Mn8@1127_g N_VSS_Mn8@1127_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1126 N_OUT8_Mn8@1126_d N_OUT7_Mn8@1126_g N_VSS_Mn8@1126_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1127 N_OUT8_Mp8@1127_d N_OUT7_Mp8@1127_g N_VDD_Mp8@1127_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1126 N_OUT8_Mp8@1126_d N_OUT7_Mp8@1126_g N_VDD_Mp8@1126_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1125 N_OUT8_Mn8@1125_d N_OUT7_Mn8@1125_g N_VSS_Mn8@1125_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1124 N_OUT8_Mn8@1124_d N_OUT7_Mn8@1124_g N_VSS_Mn8@1124_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1125 N_OUT8_Mp8@1125_d N_OUT7_Mp8@1125_g N_VDD_Mp8@1125_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1124 N_OUT8_Mp8@1124_d N_OUT7_Mp8@1124_g N_VDD_Mp8@1124_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1123 N_OUT8_Mn8@1123_d N_OUT7_Mn8@1123_g N_VSS_Mn8@1123_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1122 N_OUT8_Mn8@1122_d N_OUT7_Mn8@1122_g N_VSS_Mn8@1122_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1123 N_OUT8_Mp8@1123_d N_OUT7_Mp8@1123_g N_VDD_Mp8@1123_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1122 N_OUT8_Mp8@1122_d N_OUT7_Mp8@1122_g N_VDD_Mp8@1122_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1121 N_OUT8_Mn8@1121_d N_OUT7_Mn8@1121_g N_VSS_Mn8@1121_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1120 N_OUT8_Mn8@1120_d N_OUT7_Mn8@1120_g N_VSS_Mn8@1120_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1121 N_OUT8_Mp8@1121_d N_OUT7_Mp8@1121_g N_VDD_Mp8@1121_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1120 N_OUT8_Mp8@1120_d N_OUT7_Mp8@1120_g N_VDD_Mp8@1120_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1119 N_OUT8_Mn8@1119_d N_OUT7_Mn8@1119_g N_VSS_Mn8@1119_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1118 N_OUT8_Mn8@1118_d N_OUT7_Mn8@1118_g N_VSS_Mn8@1118_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1119 N_OUT8_Mp8@1119_d N_OUT7_Mp8@1119_g N_VDD_Mp8@1119_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1118 N_OUT8_Mp8@1118_d N_OUT7_Mp8@1118_g N_VDD_Mp8@1118_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1117 N_OUT8_Mn8@1117_d N_OUT7_Mn8@1117_g N_VSS_Mn8@1117_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1116 N_OUT8_Mn8@1116_d N_OUT7_Mn8@1116_g N_VSS_Mn8@1116_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1117 N_OUT8_Mp8@1117_d N_OUT7_Mp8@1117_g N_VDD_Mp8@1117_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1116 N_OUT8_Mp8@1116_d N_OUT7_Mp8@1116_g N_VDD_Mp8@1116_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1115 N_OUT8_Mn8@1115_d N_OUT7_Mn8@1115_g N_VSS_Mn8@1115_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1114 N_OUT8_Mn8@1114_d N_OUT7_Mn8@1114_g N_VSS_Mn8@1114_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1115 N_OUT8_Mp8@1115_d N_OUT7_Mp8@1115_g N_VDD_Mp8@1115_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1114 N_OUT8_Mp8@1114_d N_OUT7_Mp8@1114_g N_VDD_Mp8@1114_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1113 N_OUT8_Mn8@1113_d N_OUT7_Mn8@1113_g N_VSS_Mn8@1113_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1112 N_OUT8_Mn8@1112_d N_OUT7_Mn8@1112_g N_VSS_Mn8@1112_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1113 N_OUT8_Mp8@1113_d N_OUT7_Mp8@1113_g N_VDD_Mp8@1113_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1112 N_OUT8_Mp8@1112_d N_OUT7_Mp8@1112_g N_VDD_Mp8@1112_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1111 N_OUT8_Mn8@1111_d N_OUT7_Mn8@1111_g N_VSS_Mn8@1111_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1110 N_OUT8_Mn8@1110_d N_OUT7_Mn8@1110_g N_VSS_Mn8@1110_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1111 N_OUT8_Mp8@1111_d N_OUT7_Mp8@1111_g N_VDD_Mp8@1111_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1110 N_OUT8_Mp8@1110_d N_OUT7_Mp8@1110_g N_VDD_Mp8@1110_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1109 N_OUT8_Mn8@1109_d N_OUT7_Mn8@1109_g N_VSS_Mn8@1109_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1108 N_OUT8_Mn8@1108_d N_OUT7_Mn8@1108_g N_VSS_Mn8@1108_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1109 N_OUT8_Mp8@1109_d N_OUT7_Mp8@1109_g N_VDD_Mp8@1109_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1108 N_OUT8_Mp8@1108_d N_OUT7_Mp8@1108_g N_VDD_Mp8@1108_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1107 N_OUT8_Mn8@1107_d N_OUT7_Mn8@1107_g N_VSS_Mn8@1107_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1106 N_OUT8_Mn8@1106_d N_OUT7_Mn8@1106_g N_VSS_Mn8@1106_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1107 N_OUT8_Mp8@1107_d N_OUT7_Mp8@1107_g N_VDD_Mp8@1107_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1106 N_OUT8_Mp8@1106_d N_OUT7_Mp8@1106_g N_VDD_Mp8@1106_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1105 N_OUT8_Mn8@1105_d N_OUT7_Mn8@1105_g N_VSS_Mn8@1105_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1104 N_OUT8_Mn8@1104_d N_OUT7_Mn8@1104_g N_VSS_Mn8@1104_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1105 N_OUT8_Mp8@1105_d N_OUT7_Mp8@1105_g N_VDD_Mp8@1105_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1104 N_OUT8_Mp8@1104_d N_OUT7_Mp8@1104_g N_VDD_Mp8@1104_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1103 N_OUT8_Mn8@1103_d N_OUT7_Mn8@1103_g N_VSS_Mn8@1103_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1102 N_OUT8_Mn8@1102_d N_OUT7_Mn8@1102_g N_VSS_Mn8@1102_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1103 N_OUT8_Mp8@1103_d N_OUT7_Mp8@1103_g N_VDD_Mp8@1103_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1102 N_OUT8_Mp8@1102_d N_OUT7_Mp8@1102_g N_VDD_Mp8@1102_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1101 N_OUT8_Mn8@1101_d N_OUT7_Mn8@1101_g N_VSS_Mn8@1101_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1100 N_OUT8_Mn8@1100_d N_OUT7_Mn8@1100_g N_VSS_Mn8@1100_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1101 N_OUT8_Mp8@1101_d N_OUT7_Mp8@1101_g N_VDD_Mp8@1101_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1100 N_OUT8_Mp8@1100_d N_OUT7_Mp8@1100_g N_VDD_Mp8@1100_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1099 N_OUT8_Mn8@1099_d N_OUT7_Mn8@1099_g N_VSS_Mn8@1099_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1098 N_OUT8_Mn8@1098_d N_OUT7_Mn8@1098_g N_VSS_Mn8@1098_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1099 N_OUT8_Mp8@1099_d N_OUT7_Mp8@1099_g N_VDD_Mp8@1099_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1098 N_OUT8_Mp8@1098_d N_OUT7_Mp8@1098_g N_VDD_Mp8@1098_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1097 N_OUT8_Mn8@1097_d N_OUT7_Mn8@1097_g N_VSS_Mn8@1097_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1096 N_OUT8_Mn8@1096_d N_OUT7_Mn8@1096_g N_VSS_Mn8@1096_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1097 N_OUT8_Mp8@1097_d N_OUT7_Mp8@1097_g N_VDD_Mp8@1097_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1096 N_OUT8_Mp8@1096_d N_OUT7_Mp8@1096_g N_VDD_Mp8@1096_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1095 N_OUT8_Mn8@1095_d N_OUT7_Mn8@1095_g N_VSS_Mn8@1095_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1094 N_OUT8_Mn8@1094_d N_OUT7_Mn8@1094_g N_VSS_Mn8@1094_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1095 N_OUT8_Mp8@1095_d N_OUT7_Mp8@1095_g N_VDD_Mp8@1095_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1094 N_OUT8_Mp8@1094_d N_OUT7_Mp8@1094_g N_VDD_Mp8@1094_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1093 N_OUT8_Mn8@1093_d N_OUT7_Mn8@1093_g N_VSS_Mn8@1093_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1092 N_OUT8_Mn8@1092_d N_OUT7_Mn8@1092_g N_VSS_Mn8@1092_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1093 N_OUT8_Mp8@1093_d N_OUT7_Mp8@1093_g N_VDD_Mp8@1093_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1092 N_OUT8_Mp8@1092_d N_OUT7_Mp8@1092_g N_VDD_Mp8@1092_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1091 N_OUT8_Mn8@1091_d N_OUT7_Mn8@1091_g N_VSS_Mn8@1091_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1090 N_OUT8_Mn8@1090_d N_OUT7_Mn8@1090_g N_VSS_Mn8@1090_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1091 N_OUT8_Mp8@1091_d N_OUT7_Mp8@1091_g N_VDD_Mp8@1091_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1090 N_OUT8_Mp8@1090_d N_OUT7_Mp8@1090_g N_VDD_Mp8@1090_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1089 N_OUT8_Mn8@1089_d N_OUT7_Mn8@1089_g N_VSS_Mn8@1089_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1088 N_OUT8_Mn8@1088_d N_OUT7_Mn8@1088_g N_VSS_Mn8@1088_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1089 N_OUT8_Mp8@1089_d N_OUT7_Mp8@1089_g N_VDD_Mp8@1089_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1088 N_OUT8_Mp8@1088_d N_OUT7_Mp8@1088_g N_VDD_Mp8@1088_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1087 N_OUT8_Mn8@1087_d N_OUT7_Mn8@1087_g N_VSS_Mn8@1087_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1086 N_OUT8_Mn8@1086_d N_OUT7_Mn8@1086_g N_VSS_Mn8@1086_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1087 N_OUT8_Mp8@1087_d N_OUT7_Mp8@1087_g N_VDD_Mp8@1087_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1086 N_OUT8_Mp8@1086_d N_OUT7_Mp8@1086_g N_VDD_Mp8@1086_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1085 N_OUT8_Mn8@1085_d N_OUT7_Mn8@1085_g N_VSS_Mn8@1085_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1084 N_OUT8_Mn8@1084_d N_OUT7_Mn8@1084_g N_VSS_Mn8@1084_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1085 N_OUT8_Mp8@1085_d N_OUT7_Mp8@1085_g N_VDD_Mp8@1085_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1084 N_OUT8_Mp8@1084_d N_OUT7_Mp8@1084_g N_VDD_Mp8@1084_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1083 N_OUT8_Mn8@1083_d N_OUT7_Mn8@1083_g N_VSS_Mn8@1083_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1082 N_OUT8_Mn8@1082_d N_OUT7_Mn8@1082_g N_VSS_Mn8@1082_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1083 N_OUT8_Mp8@1083_d N_OUT7_Mp8@1083_g N_VDD_Mp8@1083_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1082 N_OUT8_Mp8@1082_d N_OUT7_Mp8@1082_g N_VDD_Mp8@1082_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1081 N_OUT8_Mn8@1081_d N_OUT7_Mn8@1081_g N_VSS_Mn8@1081_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1080 N_OUT8_Mn8@1080_d N_OUT7_Mn8@1080_g N_VSS_Mn8@1080_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1081 N_OUT8_Mp8@1081_d N_OUT7_Mp8@1081_g N_VDD_Mp8@1081_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1080 N_OUT8_Mp8@1080_d N_OUT7_Mp8@1080_g N_VDD_Mp8@1080_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1079 N_OUT8_Mn8@1079_d N_OUT7_Mn8@1079_g N_VSS_Mn8@1079_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1078 N_OUT8_Mn8@1078_d N_OUT7_Mn8@1078_g N_VSS_Mn8@1078_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1079 N_OUT8_Mp8@1079_d N_OUT7_Mp8@1079_g N_VDD_Mp8@1079_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1078 N_OUT8_Mp8@1078_d N_OUT7_Mp8@1078_g N_VDD_Mp8@1078_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1077 N_OUT8_Mn8@1077_d N_OUT7_Mn8@1077_g N_VSS_Mn8@1077_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1076 N_OUT8_Mn8@1076_d N_OUT7_Mn8@1076_g N_VSS_Mn8@1076_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1077 N_OUT8_Mp8@1077_d N_OUT7_Mp8@1077_g N_VDD_Mp8@1077_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1076 N_OUT8_Mp8@1076_d N_OUT7_Mp8@1076_g N_VDD_Mp8@1076_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1075 N_OUT8_Mn8@1075_d N_OUT7_Mn8@1075_g N_VSS_Mn8@1075_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1074 N_OUT8_Mn8@1074_d N_OUT7_Mn8@1074_g N_VSS_Mn8@1074_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1075 N_OUT8_Mp8@1075_d N_OUT7_Mp8@1075_g N_VDD_Mp8@1075_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1074 N_OUT8_Mp8@1074_d N_OUT7_Mp8@1074_g N_VDD_Mp8@1074_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1073 N_OUT8_Mn8@1073_d N_OUT7_Mn8@1073_g N_VSS_Mn8@1073_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1072 N_OUT8_Mn8@1072_d N_OUT7_Mn8@1072_g N_VSS_Mn8@1072_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1073 N_OUT8_Mp8@1073_d N_OUT7_Mp8@1073_g N_VDD_Mp8@1073_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1072 N_OUT8_Mp8@1072_d N_OUT7_Mp8@1072_g N_VDD_Mp8@1072_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1071 N_OUT8_Mn8@1071_d N_OUT7_Mn8@1071_g N_VSS_Mn8@1071_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1070 N_OUT8_Mn8@1070_d N_OUT7_Mn8@1070_g N_VSS_Mn8@1070_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1071 N_OUT8_Mp8@1071_d N_OUT7_Mp8@1071_g N_VDD_Mp8@1071_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1070 N_OUT8_Mp8@1070_d N_OUT7_Mp8@1070_g N_VDD_Mp8@1070_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1069 N_OUT8_Mn8@1069_d N_OUT7_Mn8@1069_g N_VSS_Mn8@1069_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1068 N_OUT8_Mn8@1068_d N_OUT7_Mn8@1068_g N_VSS_Mn8@1068_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1069 N_OUT8_Mp8@1069_d N_OUT7_Mp8@1069_g N_VDD_Mp8@1069_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1068 N_OUT8_Mp8@1068_d N_OUT7_Mp8@1068_g N_VDD_Mp8@1068_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1067 N_OUT8_Mn8@1067_d N_OUT7_Mn8@1067_g N_VSS_Mn8@1067_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1066 N_OUT8_Mn8@1066_d N_OUT7_Mn8@1066_g N_VSS_Mn8@1066_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1067 N_OUT8_Mp8@1067_d N_OUT7_Mp8@1067_g N_VDD_Mp8@1067_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1066 N_OUT8_Mp8@1066_d N_OUT7_Mp8@1066_g N_VDD_Mp8@1066_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1065 N_OUT8_Mn8@1065_d N_OUT7_Mn8@1065_g N_VSS_Mn8@1065_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1064 N_OUT8_Mn8@1064_d N_OUT7_Mn8@1064_g N_VSS_Mn8@1064_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1065 N_OUT8_Mp8@1065_d N_OUT7_Mp8@1065_g N_VDD_Mp8@1065_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1064 N_OUT8_Mp8@1064_d N_OUT7_Mp8@1064_g N_VDD_Mp8@1064_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1063 N_OUT8_Mn8@1063_d N_OUT7_Mn8@1063_g N_VSS_Mn8@1063_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1062 N_OUT8_Mn8@1062_d N_OUT7_Mn8@1062_g N_VSS_Mn8@1062_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1063 N_OUT8_Mp8@1063_d N_OUT7_Mp8@1063_g N_VDD_Mp8@1063_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1062 N_OUT8_Mp8@1062_d N_OUT7_Mp8@1062_g N_VDD_Mp8@1062_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1061 N_OUT8_Mn8@1061_d N_OUT7_Mn8@1061_g N_VSS_Mn8@1061_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1060 N_OUT8_Mn8@1060_d N_OUT7_Mn8@1060_g N_VSS_Mn8@1060_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1061 N_OUT8_Mp8@1061_d N_OUT7_Mp8@1061_g N_VDD_Mp8@1061_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1060 N_OUT8_Mp8@1060_d N_OUT7_Mp8@1060_g N_VDD_Mp8@1060_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1059 N_OUT8_Mn8@1059_d N_OUT7_Mn8@1059_g N_VSS_Mn8@1059_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1058 N_OUT8_Mn8@1058_d N_OUT7_Mn8@1058_g N_VSS_Mn8@1058_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1059 N_OUT8_Mp8@1059_d N_OUT7_Mp8@1059_g N_VDD_Mp8@1059_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1058 N_OUT8_Mp8@1058_d N_OUT7_Mp8@1058_g N_VDD_Mp8@1058_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1057 N_OUT8_Mn8@1057_d N_OUT7_Mn8@1057_g N_VSS_Mn8@1057_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1056 N_OUT8_Mn8@1056_d N_OUT7_Mn8@1056_g N_VSS_Mn8@1056_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1057 N_OUT8_Mp8@1057_d N_OUT7_Mp8@1057_g N_VDD_Mp8@1057_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1056 N_OUT8_Mp8@1056_d N_OUT7_Mp8@1056_g N_VDD_Mp8@1056_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1055 N_OUT8_Mn8@1055_d N_OUT7_Mn8@1055_g N_VSS_Mn8@1055_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1054 N_OUT8_Mn8@1054_d N_OUT7_Mn8@1054_g N_VSS_Mn8@1054_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1055 N_OUT8_Mp8@1055_d N_OUT7_Mp8@1055_g N_VDD_Mp8@1055_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1054 N_OUT8_Mp8@1054_d N_OUT7_Mp8@1054_g N_VDD_Mp8@1054_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1053 N_OUT8_Mn8@1053_d N_OUT7_Mn8@1053_g N_VSS_Mn8@1053_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1052 N_OUT8_Mn8@1052_d N_OUT7_Mn8@1052_g N_VSS_Mn8@1052_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1053 N_OUT8_Mp8@1053_d N_OUT7_Mp8@1053_g N_VDD_Mp8@1053_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1052 N_OUT8_Mp8@1052_d N_OUT7_Mp8@1052_g N_VDD_Mp8@1052_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1051 N_OUT8_Mn8@1051_d N_OUT7_Mn8@1051_g N_VSS_Mn8@1051_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1050 N_OUT8_Mn8@1050_d N_OUT7_Mn8@1050_g N_VSS_Mn8@1050_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1051 N_OUT8_Mp8@1051_d N_OUT7_Mp8@1051_g N_VDD_Mp8@1051_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1050 N_OUT8_Mp8@1050_d N_OUT7_Mp8@1050_g N_VDD_Mp8@1050_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1049 N_OUT8_Mn8@1049_d N_OUT7_Mn8@1049_g N_VSS_Mn8@1049_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1048 N_OUT8_Mn8@1048_d N_OUT7_Mn8@1048_g N_VSS_Mn8@1048_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1049 N_OUT8_Mp8@1049_d N_OUT7_Mp8@1049_g N_VDD_Mp8@1049_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1048 N_OUT8_Mp8@1048_d N_OUT7_Mp8@1048_g N_VDD_Mp8@1048_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1047 N_OUT8_Mn8@1047_d N_OUT7_Mn8@1047_g N_VSS_Mn8@1047_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1046 N_OUT8_Mn8@1046_d N_OUT7_Mn8@1046_g N_VSS_Mn8@1046_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1047 N_OUT8_Mp8@1047_d N_OUT7_Mp8@1047_g N_VDD_Mp8@1047_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1046 N_OUT8_Mp8@1046_d N_OUT7_Mp8@1046_g N_VDD_Mp8@1046_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1045 N_OUT8_Mn8@1045_d N_OUT7_Mn8@1045_g N_VSS_Mn8@1045_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1044 N_OUT8_Mn8@1044_d N_OUT7_Mn8@1044_g N_VSS_Mn8@1044_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1045 N_OUT8_Mp8@1045_d N_OUT7_Mp8@1045_g N_VDD_Mp8@1045_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1044 N_OUT8_Mp8@1044_d N_OUT7_Mp8@1044_g N_VDD_Mp8@1044_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1043 N_OUT8_Mn8@1043_d N_OUT7_Mn8@1043_g N_VSS_Mn8@1043_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1042 N_OUT8_Mn8@1042_d N_OUT7_Mn8@1042_g N_VSS_Mn8@1042_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1043 N_OUT8_Mp8@1043_d N_OUT7_Mp8@1043_g N_VDD_Mp8@1043_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1042 N_OUT8_Mp8@1042_d N_OUT7_Mp8@1042_g N_VDD_Mp8@1042_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1041 N_OUT8_Mn8@1041_d N_OUT7_Mn8@1041_g N_VSS_Mn8@1041_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1040 N_OUT8_Mn8@1040_d N_OUT7_Mn8@1040_g N_VSS_Mn8@1040_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1041 N_OUT8_Mp8@1041_d N_OUT7_Mp8@1041_g N_VDD_Mp8@1041_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1040 N_OUT8_Mp8@1040_d N_OUT7_Mp8@1040_g N_VDD_Mp8@1040_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1039 N_OUT8_Mn8@1039_d N_OUT7_Mn8@1039_g N_VSS_Mn8@1039_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1038 N_OUT8_Mn8@1038_d N_OUT7_Mn8@1038_g N_VSS_Mn8@1038_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1039 N_OUT8_Mp8@1039_d N_OUT7_Mp8@1039_g N_VDD_Mp8@1039_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1038 N_OUT8_Mp8@1038_d N_OUT7_Mp8@1038_g N_VDD_Mp8@1038_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1037 N_OUT8_Mn8@1037_d N_OUT7_Mn8@1037_g N_VSS_Mn8@1037_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1036 N_OUT8_Mn8@1036_d N_OUT7_Mn8@1036_g N_VSS_Mn8@1036_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1037 N_OUT8_Mp8@1037_d N_OUT7_Mp8@1037_g N_VDD_Mp8@1037_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1036 N_OUT8_Mp8@1036_d N_OUT7_Mp8@1036_g N_VDD_Mp8@1036_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1035 N_OUT8_Mn8@1035_d N_OUT7_Mn8@1035_g N_VSS_Mn8@1035_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1034 N_OUT8_Mn8@1034_d N_OUT7_Mn8@1034_g N_VSS_Mn8@1034_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1035 N_OUT8_Mp8@1035_d N_OUT7_Mp8@1035_g N_VDD_Mp8@1035_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1034 N_OUT8_Mp8@1034_d N_OUT7_Mp8@1034_g N_VDD_Mp8@1034_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1033 N_OUT8_Mn8@1033_d N_OUT7_Mn8@1033_g N_VSS_Mn8@1033_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1032 N_OUT8_Mn8@1032_d N_OUT7_Mn8@1032_g N_VSS_Mn8@1032_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1033 N_OUT8_Mp8@1033_d N_OUT7_Mp8@1033_g N_VDD_Mp8@1033_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1032 N_OUT8_Mp8@1032_d N_OUT7_Mp8@1032_g N_VDD_Mp8@1032_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1031 N_OUT8_Mn8@1031_d N_OUT7_Mn8@1031_g N_VSS_Mn8@1031_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1030 N_OUT8_Mn8@1030_d N_OUT7_Mn8@1030_g N_VSS_Mn8@1030_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1031 N_OUT8_Mp8@1031_d N_OUT7_Mp8@1031_g N_VDD_Mp8@1031_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1030 N_OUT8_Mp8@1030_d N_OUT7_Mp8@1030_g N_VDD_Mp8@1030_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1029 N_OUT8_Mn8@1029_d N_OUT7_Mn8@1029_g N_VSS_Mn8@1029_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1028 N_OUT8_Mn8@1028_d N_OUT7_Mn8@1028_g N_VSS_Mn8@1028_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1029 N_OUT8_Mp8@1029_d N_OUT7_Mp8@1029_g N_VDD_Mp8@1029_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1028 N_OUT8_Mp8@1028_d N_OUT7_Mp8@1028_g N_VDD_Mp8@1028_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1027 N_OUT8_Mn8@1027_d N_OUT7_Mn8@1027_g N_VSS_Mn8@1027_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1026 N_OUT8_Mn8@1026_d N_OUT7_Mn8@1026_g N_VSS_Mn8@1026_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1027 N_OUT8_Mp8@1027_d N_OUT7_Mp8@1027_g N_VDD_Mp8@1027_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1026 N_OUT8_Mp8@1026_d N_OUT7_Mp8@1026_g N_VDD_Mp8@1026_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1025 N_OUT8_Mn8@1025_d N_OUT7_Mn8@1025_g N_VSS_Mn8@1025_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1024 N_OUT8_Mn8@1024_d N_OUT7_Mn8@1024_g N_VSS_Mn8@1024_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1025 N_OUT8_Mp8@1025_d N_OUT7_Mp8@1025_g N_VDD_Mp8@1025_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1024 N_OUT8_Mp8@1024_d N_OUT7_Mp8@1024_g N_VDD_Mp8@1024_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1023 N_OUT8_Mn8@1023_d N_OUT7_Mn8@1023_g N_VSS_Mn8@1023_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1022 N_OUT8_Mn8@1022_d N_OUT7_Mn8@1022_g N_VSS_Mn8@1022_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1023 N_OUT8_Mp8@1023_d N_OUT7_Mp8@1023_g N_VDD_Mp8@1023_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1022 N_OUT8_Mp8@1022_d N_OUT7_Mp8@1022_g N_VDD_Mp8@1022_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1021 N_OUT8_Mn8@1021_d N_OUT7_Mn8@1021_g N_VSS_Mn8@1021_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1020 N_OUT8_Mn8@1020_d N_OUT7_Mn8@1020_g N_VSS_Mn8@1020_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1021 N_OUT8_Mp8@1021_d N_OUT7_Mp8@1021_g N_VDD_Mp8@1021_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1020 N_OUT8_Mp8@1020_d N_OUT7_Mp8@1020_g N_VDD_Mp8@1020_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1019 N_OUT8_Mn8@1019_d N_OUT7_Mn8@1019_g N_VSS_Mn8@1019_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1018 N_OUT8_Mn8@1018_d N_OUT7_Mn8@1018_g N_VSS_Mn8@1018_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1019 N_OUT8_Mp8@1019_d N_OUT7_Mp8@1019_g N_VDD_Mp8@1019_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1018 N_OUT8_Mp8@1018_d N_OUT7_Mp8@1018_g N_VDD_Mp8@1018_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1017 N_OUT8_Mn8@1017_d N_OUT7_Mn8@1017_g N_VSS_Mn8@1017_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1016 N_OUT8_Mn8@1016_d N_OUT7_Mn8@1016_g N_VSS_Mn8@1016_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1017 N_OUT8_Mp8@1017_d N_OUT7_Mp8@1017_g N_VDD_Mp8@1017_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1016 N_OUT8_Mp8@1016_d N_OUT7_Mp8@1016_g N_VDD_Mp8@1016_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1015 N_OUT8_Mn8@1015_d N_OUT7_Mn8@1015_g N_VSS_Mn8@1015_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1014 N_OUT8_Mn8@1014_d N_OUT7_Mn8@1014_g N_VSS_Mn8@1014_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1015 N_OUT8_Mp8@1015_d N_OUT7_Mp8@1015_g N_VDD_Mp8@1015_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1014 N_OUT8_Mp8@1014_d N_OUT7_Mp8@1014_g N_VDD_Mp8@1014_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1013 N_OUT8_Mn8@1013_d N_OUT7_Mn8@1013_g N_VSS_Mn8@1013_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1012 N_OUT8_Mn8@1012_d N_OUT7_Mn8@1012_g N_VSS_Mn8@1012_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1013 N_OUT8_Mp8@1013_d N_OUT7_Mp8@1013_g N_VDD_Mp8@1013_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1012 N_OUT8_Mp8@1012_d N_OUT7_Mp8@1012_g N_VDD_Mp8@1012_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1011 N_OUT8_Mn8@1011_d N_OUT7_Mn8@1011_g N_VSS_Mn8@1011_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1010 N_OUT8_Mn8@1010_d N_OUT7_Mn8@1010_g N_VSS_Mn8@1010_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1011 N_OUT8_Mp8@1011_d N_OUT7_Mp8@1011_g N_VDD_Mp8@1011_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1010 N_OUT8_Mp8@1010_d N_OUT7_Mp8@1010_g N_VDD_Mp8@1010_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1009 N_OUT8_Mn8@1009_d N_OUT7_Mn8@1009_g N_VSS_Mn8@1009_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1008 N_OUT8_Mn8@1008_d N_OUT7_Mn8@1008_g N_VSS_Mn8@1008_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1009 N_OUT8_Mp8@1009_d N_OUT7_Mp8@1009_g N_VDD_Mp8@1009_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1008 N_OUT8_Mp8@1008_d N_OUT7_Mp8@1008_g N_VDD_Mp8@1008_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1007 N_OUT8_Mn8@1007_d N_OUT7_Mn8@1007_g N_VSS_Mn8@1007_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1006 N_OUT8_Mn8@1006_d N_OUT7_Mn8@1006_g N_VSS_Mn8@1006_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1007 N_OUT8_Mp8@1007_d N_OUT7_Mp8@1007_g N_VDD_Mp8@1007_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1006 N_OUT8_Mp8@1006_d N_OUT7_Mp8@1006_g N_VDD_Mp8@1006_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1005 N_OUT8_Mn8@1005_d N_OUT7_Mn8@1005_g N_VSS_Mn8@1005_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1004 N_OUT8_Mn8@1004_d N_OUT7_Mn8@1004_g N_VSS_Mn8@1004_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1005 N_OUT8_Mp8@1005_d N_OUT7_Mp8@1005_g N_VDD_Mp8@1005_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1004 N_OUT8_Mp8@1004_d N_OUT7_Mp8@1004_g N_VDD_Mp8@1004_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1003 N_OUT8_Mn8@1003_d N_OUT7_Mn8@1003_g N_VSS_Mn8@1003_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1002 N_OUT8_Mn8@1002_d N_OUT7_Mn8@1002_g N_VSS_Mn8@1002_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1003 N_OUT8_Mp8@1003_d N_OUT7_Mp8@1003_g N_VDD_Mp8@1003_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1002 N_OUT8_Mp8@1002_d N_OUT7_Mp8@1002_g N_VDD_Mp8@1002_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@1001 N_OUT8_Mn8@1001_d N_OUT7_Mn8@1001_g N_VSS_Mn8@1001_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@1000 N_OUT8_Mn8@1000_d N_OUT7_Mn8@1000_g N_VSS_Mn8@1000_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@1001 N_OUT8_Mp8@1001_d N_OUT7_Mp8@1001_g N_VDD_Mp8@1001_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@1000 N_OUT8_Mp8@1000_d N_OUT7_Mp8@1000_g N_VDD_Mp8@1000_s N_VDD_Mp8@3769_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@999 N_OUT8_Mn8@999_d N_OUT7_Mn8@999_g N_VSS_Mn8@999_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@998 N_OUT8_Mn8@998_d N_OUT7_Mn8@998_g N_VSS_Mn8@998_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@999 N_OUT8_Mp8@999_d N_OUT7_Mp8@999_g N_VDD_Mp8@999_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@998 N_OUT8_Mp8@998_d N_OUT7_Mp8@998_g N_VDD_Mp8@998_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@997 N_OUT8_Mn8@997_d N_OUT7_Mn8@997_g N_VSS_Mn8@997_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@996 N_OUT8_Mn8@996_d N_OUT7_Mn8@996_g N_VSS_Mn8@996_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@997 N_OUT8_Mp8@997_d N_OUT7_Mp8@997_g N_VDD_Mp8@997_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@996 N_OUT8_Mp8@996_d N_OUT7_Mp8@996_g N_VDD_Mp8@996_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@995 N_OUT8_Mn8@995_d N_OUT7_Mn8@995_g N_VSS_Mn8@995_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@994 N_OUT8_Mn8@994_d N_OUT7_Mn8@994_g N_VSS_Mn8@994_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@995 N_OUT8_Mp8@995_d N_OUT7_Mp8@995_g N_VDD_Mp8@995_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@994 N_OUT8_Mp8@994_d N_OUT7_Mp8@994_g N_VDD_Mp8@994_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@993 N_OUT8_Mn8@993_d N_OUT7_Mn8@993_g N_VSS_Mn8@993_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@992 N_OUT8_Mn8@992_d N_OUT7_Mn8@992_g N_VSS_Mn8@992_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@993 N_OUT8_Mp8@993_d N_OUT7_Mp8@993_g N_VDD_Mp8@993_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@992 N_OUT8_Mp8@992_d N_OUT7_Mp8@992_g N_VDD_Mp8@992_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@991 N_OUT8_Mn8@991_d N_OUT7_Mn8@991_g N_VSS_Mn8@991_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@990 N_OUT8_Mn8@990_d N_OUT7_Mn8@990_g N_VSS_Mn8@990_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@991 N_OUT8_Mp8@991_d N_OUT7_Mp8@991_g N_VDD_Mp8@991_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@990 N_OUT8_Mp8@990_d N_OUT7_Mp8@990_g N_VDD_Mp8@990_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@989 N_OUT8_Mn8@989_d N_OUT7_Mn8@989_g N_VSS_Mn8@989_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@988 N_OUT8_Mn8@988_d N_OUT7_Mn8@988_g N_VSS_Mn8@988_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@989 N_OUT8_Mp8@989_d N_OUT7_Mp8@989_g N_VDD_Mp8@989_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@988 N_OUT8_Mp8@988_d N_OUT7_Mp8@988_g N_VDD_Mp8@988_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@987 N_OUT8_Mn8@987_d N_OUT7_Mn8@987_g N_VSS_Mn8@987_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@986 N_OUT8_Mn8@986_d N_OUT7_Mn8@986_g N_VSS_Mn8@986_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@987 N_OUT8_Mp8@987_d N_OUT7_Mp8@987_g N_VDD_Mp8@987_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@986 N_OUT8_Mp8@986_d N_OUT7_Mp8@986_g N_VDD_Mp8@986_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@985 N_OUT8_Mn8@985_d N_OUT7_Mn8@985_g N_VSS_Mn8@985_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@984 N_OUT8_Mn8@984_d N_OUT7_Mn8@984_g N_VSS_Mn8@984_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@985 N_OUT8_Mp8@985_d N_OUT7_Mp8@985_g N_VDD_Mp8@985_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@984 N_OUT8_Mp8@984_d N_OUT7_Mp8@984_g N_VDD_Mp8@984_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@983 N_OUT8_Mn8@983_d N_OUT7_Mn8@983_g N_VSS_Mn8@983_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@982 N_OUT8_Mn8@982_d N_OUT7_Mn8@982_g N_VSS_Mn8@982_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@983 N_OUT8_Mp8@983_d N_OUT7_Mp8@983_g N_VDD_Mp8@983_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@982 N_OUT8_Mp8@982_d N_OUT7_Mp8@982_g N_VDD_Mp8@982_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@981 N_OUT8_Mn8@981_d N_OUT7_Mn8@981_g N_VSS_Mn8@981_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@980 N_OUT8_Mn8@980_d N_OUT7_Mn8@980_g N_VSS_Mn8@980_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@981 N_OUT8_Mp8@981_d N_OUT7_Mp8@981_g N_VDD_Mp8@981_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@980 N_OUT8_Mp8@980_d N_OUT7_Mp8@980_g N_VDD_Mp8@980_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@979 N_OUT8_Mn8@979_d N_OUT7_Mn8@979_g N_VSS_Mn8@979_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@978 N_OUT8_Mn8@978_d N_OUT7_Mn8@978_g N_VSS_Mn8@978_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@979 N_OUT8_Mp8@979_d N_OUT7_Mp8@979_g N_VDD_Mp8@979_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@978 N_OUT8_Mp8@978_d N_OUT7_Mp8@978_g N_VDD_Mp8@978_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@977 N_OUT8_Mn8@977_d N_OUT7_Mn8@977_g N_VSS_Mn8@977_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@976 N_OUT8_Mn8@976_d N_OUT7_Mn8@976_g N_VSS_Mn8@976_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@977 N_OUT8_Mp8@977_d N_OUT7_Mp8@977_g N_VDD_Mp8@977_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@976 N_OUT8_Mp8@976_d N_OUT7_Mp8@976_g N_VDD_Mp8@976_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@975 N_OUT8_Mn8@975_d N_OUT7_Mn8@975_g N_VSS_Mn8@975_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@974 N_OUT8_Mn8@974_d N_OUT7_Mn8@974_g N_VSS_Mn8@974_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@975 N_OUT8_Mp8@975_d N_OUT7_Mp8@975_g N_VDD_Mp8@975_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@974 N_OUT8_Mp8@974_d N_OUT7_Mp8@974_g N_VDD_Mp8@974_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@973 N_OUT8_Mn8@973_d N_OUT7_Mn8@973_g N_VSS_Mn8@973_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@972 N_OUT8_Mn8@972_d N_OUT7_Mn8@972_g N_VSS_Mn8@972_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@973 N_OUT8_Mp8@973_d N_OUT7_Mp8@973_g N_VDD_Mp8@973_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@972 N_OUT8_Mp8@972_d N_OUT7_Mp8@972_g N_VDD_Mp8@972_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@971 N_OUT8_Mn8@971_d N_OUT7_Mn8@971_g N_VSS_Mn8@971_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@970 N_OUT8_Mn8@970_d N_OUT7_Mn8@970_g N_VSS_Mn8@970_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@971 N_OUT8_Mp8@971_d N_OUT7_Mp8@971_g N_VDD_Mp8@971_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@970 N_OUT8_Mp8@970_d N_OUT7_Mp8@970_g N_VDD_Mp8@970_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@969 N_OUT8_Mn8@969_d N_OUT7_Mn8@969_g N_VSS_Mn8@969_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@968 N_OUT8_Mn8@968_d N_OUT7_Mn8@968_g N_VSS_Mn8@968_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@969 N_OUT8_Mp8@969_d N_OUT7_Mp8@969_g N_VDD_Mp8@969_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@968 N_OUT8_Mp8@968_d N_OUT7_Mp8@968_g N_VDD_Mp8@968_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@967 N_OUT8_Mn8@967_d N_OUT7_Mn8@967_g N_VSS_Mn8@967_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@966 N_OUT8_Mn8@966_d N_OUT7_Mn8@966_g N_VSS_Mn8@966_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@967 N_OUT8_Mp8@967_d N_OUT7_Mp8@967_g N_VDD_Mp8@967_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@966 N_OUT8_Mp8@966_d N_OUT7_Mp8@966_g N_VDD_Mp8@966_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@965 N_OUT8_Mn8@965_d N_OUT7_Mn8@965_g N_VSS_Mn8@965_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@964 N_OUT8_Mn8@964_d N_OUT7_Mn8@964_g N_VSS_Mn8@964_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@965 N_OUT8_Mp8@965_d N_OUT7_Mp8@965_g N_VDD_Mp8@965_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@964 N_OUT8_Mp8@964_d N_OUT7_Mp8@964_g N_VDD_Mp8@964_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@963 N_OUT8_Mn8@963_d N_OUT7_Mn8@963_g N_VSS_Mn8@963_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@962 N_OUT8_Mn8@962_d N_OUT7_Mn8@962_g N_VSS_Mn8@962_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@963 N_OUT8_Mp8@963_d N_OUT7_Mp8@963_g N_VDD_Mp8@963_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@962 N_OUT8_Mp8@962_d N_OUT7_Mp8@962_g N_VDD_Mp8@962_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@961 N_OUT8_Mn8@961_d N_OUT7_Mn8@961_g N_VSS_Mn8@961_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@960 N_OUT8_Mn8@960_d N_OUT7_Mn8@960_g N_VSS_Mn8@960_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@961 N_OUT8_Mp8@961_d N_OUT7_Mp8@961_g N_VDD_Mp8@961_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@960 N_OUT8_Mp8@960_d N_OUT7_Mp8@960_g N_VDD_Mp8@960_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@959 N_OUT8_Mn8@959_d N_OUT7_Mn8@959_g N_VSS_Mn8@959_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@958 N_OUT8_Mn8@958_d N_OUT7_Mn8@958_g N_VSS_Mn8@958_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@959 N_OUT8_Mp8@959_d N_OUT7_Mp8@959_g N_VDD_Mp8@959_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@958 N_OUT8_Mp8@958_d N_OUT7_Mp8@958_g N_VDD_Mp8@958_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@957 N_OUT8_Mn8@957_d N_OUT7_Mn8@957_g N_VSS_Mn8@957_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@956 N_OUT8_Mn8@956_d N_OUT7_Mn8@956_g N_VSS_Mn8@956_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@957 N_OUT8_Mp8@957_d N_OUT7_Mp8@957_g N_VDD_Mp8@957_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@956 N_OUT8_Mp8@956_d N_OUT7_Mp8@956_g N_VDD_Mp8@956_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@955 N_OUT8_Mn8@955_d N_OUT7_Mn8@955_g N_VSS_Mn8@955_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@954 N_OUT8_Mn8@954_d N_OUT7_Mn8@954_g N_VSS_Mn8@954_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@955 N_OUT8_Mp8@955_d N_OUT7_Mp8@955_g N_VDD_Mp8@955_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@954 N_OUT8_Mp8@954_d N_OUT7_Mp8@954_g N_VDD_Mp8@954_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@953 N_OUT8_Mn8@953_d N_OUT7_Mn8@953_g N_VSS_Mn8@953_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@952 N_OUT8_Mn8@952_d N_OUT7_Mn8@952_g N_VSS_Mn8@952_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@953 N_OUT8_Mp8@953_d N_OUT7_Mp8@953_g N_VDD_Mp8@953_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@952 N_OUT8_Mp8@952_d N_OUT7_Mp8@952_g N_VDD_Mp8@952_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@951 N_OUT8_Mn8@951_d N_OUT7_Mn8@951_g N_VSS_Mn8@951_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@950 N_OUT8_Mn8@950_d N_OUT7_Mn8@950_g N_VSS_Mn8@950_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@951 N_OUT8_Mp8@951_d N_OUT7_Mp8@951_g N_VDD_Mp8@951_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@950 N_OUT8_Mp8@950_d N_OUT7_Mp8@950_g N_VDD_Mp8@950_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@949 N_OUT8_Mn8@949_d N_OUT7_Mn8@949_g N_VSS_Mn8@949_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@948 N_OUT8_Mn8@948_d N_OUT7_Mn8@948_g N_VSS_Mn8@948_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@949 N_OUT8_Mp8@949_d N_OUT7_Mp8@949_g N_VDD_Mp8@949_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@948 N_OUT8_Mp8@948_d N_OUT7_Mp8@948_g N_VDD_Mp8@948_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@947 N_OUT8_Mn8@947_d N_OUT7_Mn8@947_g N_VSS_Mn8@947_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@946 N_OUT8_Mn8@946_d N_OUT7_Mn8@946_g N_VSS_Mn8@946_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@947 N_OUT8_Mp8@947_d N_OUT7_Mp8@947_g N_VDD_Mp8@947_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@946 N_OUT8_Mp8@946_d N_OUT7_Mp8@946_g N_VDD_Mp8@946_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@945 N_OUT8_Mn8@945_d N_OUT7_Mn8@945_g N_VSS_Mn8@945_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@944 N_OUT8_Mn8@944_d N_OUT7_Mn8@944_g N_VSS_Mn8@944_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@945 N_OUT8_Mp8@945_d N_OUT7_Mp8@945_g N_VDD_Mp8@945_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@944 N_OUT8_Mp8@944_d N_OUT7_Mp8@944_g N_VDD_Mp8@944_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@943 N_OUT8_Mn8@943_d N_OUT7_Mn8@943_g N_VSS_Mn8@943_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@942 N_OUT8_Mn8@942_d N_OUT7_Mn8@942_g N_VSS_Mn8@942_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@943 N_OUT8_Mp8@943_d N_OUT7_Mp8@943_g N_VDD_Mp8@943_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@942 N_OUT8_Mp8@942_d N_OUT7_Mp8@942_g N_VDD_Mp8@942_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@941 N_OUT8_Mn8@941_d N_OUT7_Mn8@941_g N_VSS_Mn8@941_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@940 N_OUT8_Mn8@940_d N_OUT7_Mn8@940_g N_VSS_Mn8@940_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@941 N_OUT8_Mp8@941_d N_OUT7_Mp8@941_g N_VDD_Mp8@941_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@940 N_OUT8_Mp8@940_d N_OUT7_Mp8@940_g N_VDD_Mp8@940_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@939 N_OUT8_Mn8@939_d N_OUT7_Mn8@939_g N_VSS_Mn8@939_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@938 N_OUT8_Mn8@938_d N_OUT7_Mn8@938_g N_VSS_Mn8@938_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@939 N_OUT8_Mp8@939_d N_OUT7_Mp8@939_g N_VDD_Mp8@939_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@938 N_OUT8_Mp8@938_d N_OUT7_Mp8@938_g N_VDD_Mp8@938_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@937 N_OUT8_Mn8@937_d N_OUT7_Mn8@937_g N_VSS_Mn8@937_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@936 N_OUT8_Mn8@936_d N_OUT7_Mn8@936_g N_VSS_Mn8@936_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@937 N_OUT8_Mp8@937_d N_OUT7_Mp8@937_g N_VDD_Mp8@937_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@936 N_OUT8_Mp8@936_d N_OUT7_Mp8@936_g N_VDD_Mp8@936_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@935 N_OUT8_Mn8@935_d N_OUT7_Mn8@935_g N_VSS_Mn8@935_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@934 N_OUT8_Mn8@934_d N_OUT7_Mn8@934_g N_VSS_Mn8@934_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@935 N_OUT8_Mp8@935_d N_OUT7_Mp8@935_g N_VDD_Mp8@935_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@934 N_OUT8_Mp8@934_d N_OUT7_Mp8@934_g N_VDD_Mp8@934_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@933 N_OUT8_Mn8@933_d N_OUT7_Mn8@933_g N_VSS_Mn8@933_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@932 N_OUT8_Mn8@932_d N_OUT7_Mn8@932_g N_VSS_Mn8@932_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@933 N_OUT8_Mp8@933_d N_OUT7_Mp8@933_g N_VDD_Mp8@933_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@932 N_OUT8_Mp8@932_d N_OUT7_Mp8@932_g N_VDD_Mp8@932_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@931 N_OUT8_Mn8@931_d N_OUT7_Mn8@931_g N_VSS_Mn8@931_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@930 N_OUT8_Mn8@930_d N_OUT7_Mn8@930_g N_VSS_Mn8@930_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@931 N_OUT8_Mp8@931_d N_OUT7_Mp8@931_g N_VDD_Mp8@931_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@930 N_OUT8_Mp8@930_d N_OUT7_Mp8@930_g N_VDD_Mp8@930_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@929 N_OUT8_Mn8@929_d N_OUT7_Mn8@929_g N_VSS_Mn8@929_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@928 N_OUT8_Mn8@928_d N_OUT7_Mn8@928_g N_VSS_Mn8@928_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@929 N_OUT8_Mp8@929_d N_OUT7_Mp8@929_g N_VDD_Mp8@929_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@928 N_OUT8_Mp8@928_d N_OUT7_Mp8@928_g N_VDD_Mp8@928_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@927 N_OUT8_Mn8@927_d N_OUT7_Mn8@927_g N_VSS_Mn8@927_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@926 N_OUT8_Mn8@926_d N_OUT7_Mn8@926_g N_VSS_Mn8@926_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@927 N_OUT8_Mp8@927_d N_OUT7_Mp8@927_g N_VDD_Mp8@927_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@926 N_OUT8_Mp8@926_d N_OUT7_Mp8@926_g N_VDD_Mp8@926_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@925 N_OUT8_Mn8@925_d N_OUT7_Mn8@925_g N_VSS_Mn8@925_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@924 N_OUT8_Mn8@924_d N_OUT7_Mn8@924_g N_VSS_Mn8@924_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@925 N_OUT8_Mp8@925_d N_OUT7_Mp8@925_g N_VDD_Mp8@925_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@924 N_OUT8_Mp8@924_d N_OUT7_Mp8@924_g N_VDD_Mp8@924_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@923 N_OUT8_Mn8@923_d N_OUT7_Mn8@923_g N_VSS_Mn8@923_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@922 N_OUT8_Mn8@922_d N_OUT7_Mn8@922_g N_VSS_Mn8@922_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@923 N_OUT8_Mp8@923_d N_OUT7_Mp8@923_g N_VDD_Mp8@923_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@922 N_OUT8_Mp8@922_d N_OUT7_Mp8@922_g N_VDD_Mp8@922_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@921 N_OUT8_Mn8@921_d N_OUT7_Mn8@921_g N_VSS_Mn8@921_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@920 N_OUT8_Mn8@920_d N_OUT7_Mn8@920_g N_VSS_Mn8@920_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@921 N_OUT8_Mp8@921_d N_OUT7_Mp8@921_g N_VDD_Mp8@921_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@920 N_OUT8_Mp8@920_d N_OUT7_Mp8@920_g N_VDD_Mp8@920_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@919 N_OUT8_Mn8@919_d N_OUT7_Mn8@919_g N_VSS_Mn8@919_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@918 N_OUT8_Mn8@918_d N_OUT7_Mn8@918_g N_VSS_Mn8@918_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@919 N_OUT8_Mp8@919_d N_OUT7_Mp8@919_g N_VDD_Mp8@919_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@918 N_OUT8_Mp8@918_d N_OUT7_Mp8@918_g N_VDD_Mp8@918_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@917 N_OUT8_Mn8@917_d N_OUT7_Mn8@917_g N_VSS_Mn8@917_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@916 N_OUT8_Mn8@916_d N_OUT7_Mn8@916_g N_VSS_Mn8@916_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@917 N_OUT8_Mp8@917_d N_OUT7_Mp8@917_g N_VDD_Mp8@917_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@916 N_OUT8_Mp8@916_d N_OUT7_Mp8@916_g N_VDD_Mp8@916_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@915 N_OUT8_Mn8@915_d N_OUT7_Mn8@915_g N_VSS_Mn8@915_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@914 N_OUT8_Mn8@914_d N_OUT7_Mn8@914_g N_VSS_Mn8@914_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@915 N_OUT8_Mp8@915_d N_OUT7_Mp8@915_g N_VDD_Mp8@915_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@914 N_OUT8_Mp8@914_d N_OUT7_Mp8@914_g N_VDD_Mp8@914_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@913 N_OUT8_Mn8@913_d N_OUT7_Mn8@913_g N_VSS_Mn8@913_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@912 N_OUT8_Mn8@912_d N_OUT7_Mn8@912_g N_VSS_Mn8@912_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@913 N_OUT8_Mp8@913_d N_OUT7_Mp8@913_g N_VDD_Mp8@913_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@912 N_OUT8_Mp8@912_d N_OUT7_Mp8@912_g N_VDD_Mp8@912_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@911 N_OUT8_Mn8@911_d N_OUT7_Mn8@911_g N_VSS_Mn8@911_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@910 N_OUT8_Mn8@910_d N_OUT7_Mn8@910_g N_VSS_Mn8@910_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@911 N_OUT8_Mp8@911_d N_OUT7_Mp8@911_g N_VDD_Mp8@911_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@910 N_OUT8_Mp8@910_d N_OUT7_Mp8@910_g N_VDD_Mp8@910_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@909 N_OUT8_Mn8@909_d N_OUT7_Mn8@909_g N_VSS_Mn8@909_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@908 N_OUT8_Mn8@908_d N_OUT7_Mn8@908_g N_VSS_Mn8@908_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@909 N_OUT8_Mp8@909_d N_OUT7_Mp8@909_g N_VDD_Mp8@909_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@908 N_OUT8_Mp8@908_d N_OUT7_Mp8@908_g N_VDD_Mp8@908_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@907 N_OUT8_Mn8@907_d N_OUT7_Mn8@907_g N_VSS_Mn8@907_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@906 N_OUT8_Mn8@906_d N_OUT7_Mn8@906_g N_VSS_Mn8@906_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@907 N_OUT8_Mp8@907_d N_OUT7_Mp8@907_g N_VDD_Mp8@907_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@906 N_OUT8_Mp8@906_d N_OUT7_Mp8@906_g N_VDD_Mp8@906_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@905 N_OUT8_Mn8@905_d N_OUT7_Mn8@905_g N_VSS_Mn8@905_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@904 N_OUT8_Mn8@904_d N_OUT7_Mn8@904_g N_VSS_Mn8@904_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@905 N_OUT8_Mp8@905_d N_OUT7_Mp8@905_g N_VDD_Mp8@905_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@904 N_OUT8_Mp8@904_d N_OUT7_Mp8@904_g N_VDD_Mp8@904_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@903 N_OUT8_Mn8@903_d N_OUT7_Mn8@903_g N_VSS_Mn8@903_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@902 N_OUT8_Mn8@902_d N_OUT7_Mn8@902_g N_VSS_Mn8@902_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@903 N_OUT8_Mp8@903_d N_OUT7_Mp8@903_g N_VDD_Mp8@903_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@902 N_OUT8_Mp8@902_d N_OUT7_Mp8@902_g N_VDD_Mp8@902_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@901 N_OUT8_Mn8@901_d N_OUT7_Mn8@901_g N_VSS_Mn8@901_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@900 N_OUT8_Mn8@900_d N_OUT7_Mn8@900_g N_VSS_Mn8@900_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@901 N_OUT8_Mp8@901_d N_OUT7_Mp8@901_g N_VDD_Mp8@901_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@900 N_OUT8_Mp8@900_d N_OUT7_Mp8@900_g N_VDD_Mp8@900_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@899 N_OUT8_Mn8@899_d N_OUT7_Mn8@899_g N_VSS_Mn8@899_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@898 N_OUT8_Mn8@898_d N_OUT7_Mn8@898_g N_VSS_Mn8@898_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@899 N_OUT8_Mp8@899_d N_OUT7_Mp8@899_g N_VDD_Mp8@899_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@898 N_OUT8_Mp8@898_d N_OUT7_Mp8@898_g N_VDD_Mp8@898_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@897 N_OUT8_Mn8@897_d N_OUT7_Mn8@897_g N_VSS_Mn8@897_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@896 N_OUT8_Mn8@896_d N_OUT7_Mn8@896_g N_VSS_Mn8@896_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@897 N_OUT8_Mp8@897_d N_OUT7_Mp8@897_g N_VDD_Mp8@897_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@896 N_OUT8_Mp8@896_d N_OUT7_Mp8@896_g N_VDD_Mp8@896_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@895 N_OUT8_Mn8@895_d N_OUT7_Mn8@895_g N_VSS_Mn8@895_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@894 N_OUT8_Mn8@894_d N_OUT7_Mn8@894_g N_VSS_Mn8@894_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@895 N_OUT8_Mp8@895_d N_OUT7_Mp8@895_g N_VDD_Mp8@895_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@894 N_OUT8_Mp8@894_d N_OUT7_Mp8@894_g N_VDD_Mp8@894_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@893 N_OUT8_Mn8@893_d N_OUT7_Mn8@893_g N_VSS_Mn8@893_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@892 N_OUT8_Mn8@892_d N_OUT7_Mn8@892_g N_VSS_Mn8@892_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@893 N_OUT8_Mp8@893_d N_OUT7_Mp8@893_g N_VDD_Mp8@893_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@892 N_OUT8_Mp8@892_d N_OUT7_Mp8@892_g N_VDD_Mp8@892_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@891 N_OUT8_Mn8@891_d N_OUT7_Mn8@891_g N_VSS_Mn8@891_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@890 N_OUT8_Mn8@890_d N_OUT7_Mn8@890_g N_VSS_Mn8@890_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@891 N_OUT8_Mp8@891_d N_OUT7_Mp8@891_g N_VDD_Mp8@891_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@890 N_OUT8_Mp8@890_d N_OUT7_Mp8@890_g N_VDD_Mp8@890_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@889 N_OUT8_Mn8@889_d N_OUT7_Mn8@889_g N_VSS_Mn8@889_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@888 N_OUT8_Mn8@888_d N_OUT7_Mn8@888_g N_VSS_Mn8@888_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@889 N_OUT8_Mp8@889_d N_OUT7_Mp8@889_g N_VDD_Mp8@889_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@888 N_OUT8_Mp8@888_d N_OUT7_Mp8@888_g N_VDD_Mp8@888_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@887 N_OUT8_Mn8@887_d N_OUT7_Mn8@887_g N_VSS_Mn8@887_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@886 N_OUT8_Mn8@886_d N_OUT7_Mn8@886_g N_VSS_Mn8@886_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@887 N_OUT8_Mp8@887_d N_OUT7_Mp8@887_g N_VDD_Mp8@887_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@886 N_OUT8_Mp8@886_d N_OUT7_Mp8@886_g N_VDD_Mp8@886_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@885 N_OUT8_Mn8@885_d N_OUT7_Mn8@885_g N_VSS_Mn8@885_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@884 N_OUT8_Mn8@884_d N_OUT7_Mn8@884_g N_VSS_Mn8@884_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@885 N_OUT8_Mp8@885_d N_OUT7_Mp8@885_g N_VDD_Mp8@885_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@884 N_OUT8_Mp8@884_d N_OUT7_Mp8@884_g N_VDD_Mp8@884_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@883 N_OUT8_Mn8@883_d N_OUT7_Mn8@883_g N_VSS_Mn8@883_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@882 N_OUT8_Mn8@882_d N_OUT7_Mn8@882_g N_VSS_Mn8@882_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@883 N_OUT8_Mp8@883_d N_OUT7_Mp8@883_g N_VDD_Mp8@883_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@882 N_OUT8_Mp8@882_d N_OUT7_Mp8@882_g N_VDD_Mp8@882_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@881 N_OUT8_Mn8@881_d N_OUT7_Mn8@881_g N_VSS_Mn8@881_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@880 N_OUT8_Mn8@880_d N_OUT7_Mn8@880_g N_VSS_Mn8@880_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@881 N_OUT8_Mp8@881_d N_OUT7_Mp8@881_g N_VDD_Mp8@881_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@880 N_OUT8_Mp8@880_d N_OUT7_Mp8@880_g N_VDD_Mp8@880_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@879 N_OUT8_Mn8@879_d N_OUT7_Mn8@879_g N_VSS_Mn8@879_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@878 N_OUT8_Mn8@878_d N_OUT7_Mn8@878_g N_VSS_Mn8@878_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@879 N_OUT8_Mp8@879_d N_OUT7_Mp8@879_g N_VDD_Mp8@879_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@878 N_OUT8_Mp8@878_d N_OUT7_Mp8@878_g N_VDD_Mp8@878_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@877 N_OUT8_Mn8@877_d N_OUT7_Mn8@877_g N_VSS_Mn8@877_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@876 N_OUT8_Mn8@876_d N_OUT7_Mn8@876_g N_VSS_Mn8@876_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@877 N_OUT8_Mp8@877_d N_OUT7_Mp8@877_g N_VDD_Mp8@877_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@876 N_OUT8_Mp8@876_d N_OUT7_Mp8@876_g N_VDD_Mp8@876_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@875 N_OUT8_Mn8@875_d N_OUT7_Mn8@875_g N_VSS_Mn8@875_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@874 N_OUT8_Mn8@874_d N_OUT7_Mn8@874_g N_VSS_Mn8@874_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@875 N_OUT8_Mp8@875_d N_OUT7_Mp8@875_g N_VDD_Mp8@875_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@874 N_OUT8_Mp8@874_d N_OUT7_Mp8@874_g N_VDD_Mp8@874_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@873 N_OUT8_Mn8@873_d N_OUT7_Mn8@873_g N_VSS_Mn8@873_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@872 N_OUT8_Mn8@872_d N_OUT7_Mn8@872_g N_VSS_Mn8@872_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@873 N_OUT8_Mp8@873_d N_OUT7_Mp8@873_g N_VDD_Mp8@873_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@872 N_OUT8_Mp8@872_d N_OUT7_Mp8@872_g N_VDD_Mp8@872_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@871 N_OUT8_Mn8@871_d N_OUT7_Mn8@871_g N_VSS_Mn8@871_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@870 N_OUT8_Mn8@870_d N_OUT7_Mn8@870_g N_VSS_Mn8@870_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@871 N_OUT8_Mp8@871_d N_OUT7_Mp8@871_g N_VDD_Mp8@871_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@870 N_OUT8_Mp8@870_d N_OUT7_Mp8@870_g N_VDD_Mp8@870_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@869 N_OUT8_Mn8@869_d N_OUT7_Mn8@869_g N_VSS_Mn8@869_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@868 N_OUT8_Mn8@868_d N_OUT7_Mn8@868_g N_VSS_Mn8@868_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@869 N_OUT8_Mp8@869_d N_OUT7_Mp8@869_g N_VDD_Mp8@869_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@868 N_OUT8_Mp8@868_d N_OUT7_Mp8@868_g N_VDD_Mp8@868_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@867 N_OUT8_Mn8@867_d N_OUT7_Mn8@867_g N_VSS_Mn8@867_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@866 N_OUT8_Mn8@866_d N_OUT7_Mn8@866_g N_VSS_Mn8@866_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@867 N_OUT8_Mp8@867_d N_OUT7_Mp8@867_g N_VDD_Mp8@867_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@866 N_OUT8_Mp8@866_d N_OUT7_Mp8@866_g N_VDD_Mp8@866_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@865 N_OUT8_Mn8@865_d N_OUT7_Mn8@865_g N_VSS_Mn8@865_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@864 N_OUT8_Mn8@864_d N_OUT7_Mn8@864_g N_VSS_Mn8@864_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@865 N_OUT8_Mp8@865_d N_OUT7_Mp8@865_g N_VDD_Mp8@865_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@864 N_OUT8_Mp8@864_d N_OUT7_Mp8@864_g N_VDD_Mp8@864_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@863 N_OUT8_Mn8@863_d N_OUT7_Mn8@863_g N_VSS_Mn8@863_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@862 N_OUT8_Mn8@862_d N_OUT7_Mn8@862_g N_VSS_Mn8@862_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@863 N_OUT8_Mp8@863_d N_OUT7_Mp8@863_g N_VDD_Mp8@863_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@862 N_OUT8_Mp8@862_d N_OUT7_Mp8@862_g N_VDD_Mp8@862_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@861 N_OUT8_Mn8@861_d N_OUT7_Mn8@861_g N_VSS_Mn8@861_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@860 N_OUT8_Mn8@860_d N_OUT7_Mn8@860_g N_VSS_Mn8@860_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@861 N_OUT8_Mp8@861_d N_OUT7_Mp8@861_g N_VDD_Mp8@861_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@860 N_OUT8_Mp8@860_d N_OUT7_Mp8@860_g N_VDD_Mp8@860_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@859 N_OUT8_Mn8@859_d N_OUT7_Mn8@859_g N_VSS_Mn8@859_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@858 N_OUT8_Mn8@858_d N_OUT7_Mn8@858_g N_VSS_Mn8@858_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@859 N_OUT8_Mp8@859_d N_OUT7_Mp8@859_g N_VDD_Mp8@859_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@858 N_OUT8_Mp8@858_d N_OUT7_Mp8@858_g N_VDD_Mp8@858_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@857 N_OUT8_Mn8@857_d N_OUT7_Mn8@857_g N_VSS_Mn8@857_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@856 N_OUT8_Mn8@856_d N_OUT7_Mn8@856_g N_VSS_Mn8@856_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@857 N_OUT8_Mp8@857_d N_OUT7_Mp8@857_g N_VDD_Mp8@857_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@856 N_OUT8_Mp8@856_d N_OUT7_Mp8@856_g N_VDD_Mp8@856_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@855 N_OUT8_Mn8@855_d N_OUT7_Mn8@855_g N_VSS_Mn8@855_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@854 N_OUT8_Mn8@854_d N_OUT7_Mn8@854_g N_VSS_Mn8@854_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@855 N_OUT8_Mp8@855_d N_OUT7_Mp8@855_g N_VDD_Mp8@855_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@854 N_OUT8_Mp8@854_d N_OUT7_Mp8@854_g N_VDD_Mp8@854_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@853 N_OUT8_Mn8@853_d N_OUT7_Mn8@853_g N_VSS_Mn8@853_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@852 N_OUT8_Mn8@852_d N_OUT7_Mn8@852_g N_VSS_Mn8@852_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@853 N_OUT8_Mp8@853_d N_OUT7_Mp8@853_g N_VDD_Mp8@853_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@852 N_OUT8_Mp8@852_d N_OUT7_Mp8@852_g N_VDD_Mp8@852_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@851 N_OUT8_Mn8@851_d N_OUT7_Mn8@851_g N_VSS_Mn8@851_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@850 N_OUT8_Mn8@850_d N_OUT7_Mn8@850_g N_VSS_Mn8@850_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@851 N_OUT8_Mp8@851_d N_OUT7_Mp8@851_g N_VDD_Mp8@851_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@850 N_OUT8_Mp8@850_d N_OUT7_Mp8@850_g N_VDD_Mp8@850_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@849 N_OUT8_Mn8@849_d N_OUT7_Mn8@849_g N_VSS_Mn8@849_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@848 N_OUT8_Mn8@848_d N_OUT7_Mn8@848_g N_VSS_Mn8@848_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@849 N_OUT8_Mp8@849_d N_OUT7_Mp8@849_g N_VDD_Mp8@849_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@848 N_OUT8_Mp8@848_d N_OUT7_Mp8@848_g N_VDD_Mp8@848_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@847 N_OUT8_Mn8@847_d N_OUT7_Mn8@847_g N_VSS_Mn8@847_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@846 N_OUT8_Mn8@846_d N_OUT7_Mn8@846_g N_VSS_Mn8@846_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@847 N_OUT8_Mp8@847_d N_OUT7_Mp8@847_g N_VDD_Mp8@847_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@846 N_OUT8_Mp8@846_d N_OUT7_Mp8@846_g N_VDD_Mp8@846_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@845 N_OUT8_Mn8@845_d N_OUT7_Mn8@845_g N_VSS_Mn8@845_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@844 N_OUT8_Mn8@844_d N_OUT7_Mn8@844_g N_VSS_Mn8@844_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@845 N_OUT8_Mp8@845_d N_OUT7_Mp8@845_g N_VDD_Mp8@845_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@844 N_OUT8_Mp8@844_d N_OUT7_Mp8@844_g N_VDD_Mp8@844_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@843 N_OUT8_Mn8@843_d N_OUT7_Mn8@843_g N_VSS_Mn8@843_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@842 N_OUT8_Mn8@842_d N_OUT7_Mn8@842_g N_VSS_Mn8@842_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@843 N_OUT8_Mp8@843_d N_OUT7_Mp8@843_g N_VDD_Mp8@843_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@842 N_OUT8_Mp8@842_d N_OUT7_Mp8@842_g N_VDD_Mp8@842_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@841 N_OUT8_Mn8@841_d N_OUT7_Mn8@841_g N_VSS_Mn8@841_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@840 N_OUT8_Mn8@840_d N_OUT7_Mn8@840_g N_VSS_Mn8@840_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@841 N_OUT8_Mp8@841_d N_OUT7_Mp8@841_g N_VDD_Mp8@841_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@840 N_OUT8_Mp8@840_d N_OUT7_Mp8@840_g N_VDD_Mp8@840_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@839 N_OUT8_Mn8@839_d N_OUT7_Mn8@839_g N_VSS_Mn8@839_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@838 N_OUT8_Mn8@838_d N_OUT7_Mn8@838_g N_VSS_Mn8@838_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@839 N_OUT8_Mp8@839_d N_OUT7_Mp8@839_g N_VDD_Mp8@839_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@838 N_OUT8_Mp8@838_d N_OUT7_Mp8@838_g N_VDD_Mp8@838_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@837 N_OUT8_Mn8@837_d N_OUT7_Mn8@837_g N_VSS_Mn8@837_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@836 N_OUT8_Mn8@836_d N_OUT7_Mn8@836_g N_VSS_Mn8@836_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@837 N_OUT8_Mp8@837_d N_OUT7_Mp8@837_g N_VDD_Mp8@837_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@836 N_OUT8_Mp8@836_d N_OUT7_Mp8@836_g N_VDD_Mp8@836_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@835 N_OUT8_Mn8@835_d N_OUT7_Mn8@835_g N_VSS_Mn8@835_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@834 N_OUT8_Mn8@834_d N_OUT7_Mn8@834_g N_VSS_Mn8@834_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@835 N_OUT8_Mp8@835_d N_OUT7_Mp8@835_g N_VDD_Mp8@835_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@834 N_OUT8_Mp8@834_d N_OUT7_Mp8@834_g N_VDD_Mp8@834_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@833 N_OUT8_Mn8@833_d N_OUT7_Mn8@833_g N_VSS_Mn8@833_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@832 N_OUT8_Mn8@832_d N_OUT7_Mn8@832_g N_VSS_Mn8@832_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@833 N_OUT8_Mp8@833_d N_OUT7_Mp8@833_g N_VDD_Mp8@833_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@832 N_OUT8_Mp8@832_d N_OUT7_Mp8@832_g N_VDD_Mp8@832_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@831 N_OUT8_Mn8@831_d N_OUT7_Mn8@831_g N_VSS_Mn8@831_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@830 N_OUT8_Mn8@830_d N_OUT7_Mn8@830_g N_VSS_Mn8@830_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@831 N_OUT8_Mp8@831_d N_OUT7_Mp8@831_g N_VDD_Mp8@831_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@830 N_OUT8_Mp8@830_d N_OUT7_Mp8@830_g N_VDD_Mp8@830_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@829 N_OUT8_Mn8@829_d N_OUT7_Mn8@829_g N_VSS_Mn8@829_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@828 N_OUT8_Mn8@828_d N_OUT7_Mn8@828_g N_VSS_Mn8@828_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@829 N_OUT8_Mp8@829_d N_OUT7_Mp8@829_g N_VDD_Mp8@829_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@828 N_OUT8_Mp8@828_d N_OUT7_Mp8@828_g N_VDD_Mp8@828_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@827 N_OUT8_Mn8@827_d N_OUT7_Mn8@827_g N_VSS_Mn8@827_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@826 N_OUT8_Mn8@826_d N_OUT7_Mn8@826_g N_VSS_Mn8@826_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@827 N_OUT8_Mp8@827_d N_OUT7_Mp8@827_g N_VDD_Mp8@827_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@826 N_OUT8_Mp8@826_d N_OUT7_Mp8@826_g N_VDD_Mp8@826_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@825 N_OUT8_Mn8@825_d N_OUT7_Mn8@825_g N_VSS_Mn8@825_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@824 N_OUT8_Mn8@824_d N_OUT7_Mn8@824_g N_VSS_Mn8@824_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@825 N_OUT8_Mp8@825_d N_OUT7_Mp8@825_g N_VDD_Mp8@825_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@824 N_OUT8_Mp8@824_d N_OUT7_Mp8@824_g N_VDD_Mp8@824_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@823 N_OUT8_Mn8@823_d N_OUT7_Mn8@823_g N_VSS_Mn8@823_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@822 N_OUT8_Mn8@822_d N_OUT7_Mn8@822_g N_VSS_Mn8@822_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@823 N_OUT8_Mp8@823_d N_OUT7_Mp8@823_g N_VDD_Mp8@823_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@822 N_OUT8_Mp8@822_d N_OUT7_Mp8@822_g N_VDD_Mp8@822_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@821 N_OUT8_Mn8@821_d N_OUT7_Mn8@821_g N_VSS_Mn8@821_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@820 N_OUT8_Mn8@820_d N_OUT7_Mn8@820_g N_VSS_Mn8@820_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@821 N_OUT8_Mp8@821_d N_OUT7_Mp8@821_g N_VDD_Mp8@821_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@820 N_OUT8_Mp8@820_d N_OUT7_Mp8@820_g N_VDD_Mp8@820_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@819 N_OUT8_Mn8@819_d N_OUT7_Mn8@819_g N_VSS_Mn8@819_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@818 N_OUT8_Mn8@818_d N_OUT7_Mn8@818_g N_VSS_Mn8@818_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@819 N_OUT8_Mp8@819_d N_OUT7_Mp8@819_g N_VDD_Mp8@819_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@818 N_OUT8_Mp8@818_d N_OUT7_Mp8@818_g N_VDD_Mp8@818_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@817 N_OUT8_Mn8@817_d N_OUT7_Mn8@817_g N_VSS_Mn8@817_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@816 N_OUT8_Mn8@816_d N_OUT7_Mn8@816_g N_VSS_Mn8@816_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@817 N_OUT8_Mp8@817_d N_OUT7_Mp8@817_g N_VDD_Mp8@817_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@816 N_OUT8_Mp8@816_d N_OUT7_Mp8@816_g N_VDD_Mp8@816_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@815 N_OUT8_Mn8@815_d N_OUT7_Mn8@815_g N_VSS_Mn8@815_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@814 N_OUT8_Mn8@814_d N_OUT7_Mn8@814_g N_VSS_Mn8@814_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@815 N_OUT8_Mp8@815_d N_OUT7_Mp8@815_g N_VDD_Mp8@815_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@814 N_OUT8_Mp8@814_d N_OUT7_Mp8@814_g N_VDD_Mp8@814_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@813 N_OUT8_Mn8@813_d N_OUT7_Mn8@813_g N_VSS_Mn8@813_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@812 N_OUT8_Mn8@812_d N_OUT7_Mn8@812_g N_VSS_Mn8@812_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@813 N_OUT8_Mp8@813_d N_OUT7_Mp8@813_g N_VDD_Mp8@813_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@812 N_OUT8_Mp8@812_d N_OUT7_Mp8@812_g N_VDD_Mp8@812_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@811 N_OUT8_Mn8@811_d N_OUT7_Mn8@811_g N_VSS_Mn8@811_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@810 N_OUT8_Mn8@810_d N_OUT7_Mn8@810_g N_VSS_Mn8@810_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@811 N_OUT8_Mp8@811_d N_OUT7_Mp8@811_g N_VDD_Mp8@811_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@810 N_OUT8_Mp8@810_d N_OUT7_Mp8@810_g N_VDD_Mp8@810_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@809 N_OUT8_Mn8@809_d N_OUT7_Mn8@809_g N_VSS_Mn8@809_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@808 N_OUT8_Mn8@808_d N_OUT7_Mn8@808_g N_VSS_Mn8@808_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@809 N_OUT8_Mp8@809_d N_OUT7_Mp8@809_g N_VDD_Mp8@809_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@808 N_OUT8_Mp8@808_d N_OUT7_Mp8@808_g N_VDD_Mp8@808_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@807 N_OUT8_Mn8@807_d N_OUT7_Mn8@807_g N_VSS_Mn8@807_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@806 N_OUT8_Mn8@806_d N_OUT7_Mn8@806_g N_VSS_Mn8@806_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@807 N_OUT8_Mp8@807_d N_OUT7_Mp8@807_g N_VDD_Mp8@807_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@806 N_OUT8_Mp8@806_d N_OUT7_Mp8@806_g N_VDD_Mp8@806_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@805 N_OUT8_Mn8@805_d N_OUT7_Mn8@805_g N_VSS_Mn8@805_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@804 N_OUT8_Mn8@804_d N_OUT7_Mn8@804_g N_VSS_Mn8@804_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@805 N_OUT8_Mp8@805_d N_OUT7_Mp8@805_g N_VDD_Mp8@805_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@804 N_OUT8_Mp8@804_d N_OUT7_Mp8@804_g N_VDD_Mp8@804_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@803 N_OUT8_Mn8@803_d N_OUT7_Mn8@803_g N_VSS_Mn8@803_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@802 N_OUT8_Mn8@802_d N_OUT7_Mn8@802_g N_VSS_Mn8@802_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@803 N_OUT8_Mp8@803_d N_OUT7_Mp8@803_g N_VDD_Mp8@803_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@802 N_OUT8_Mp8@802_d N_OUT7_Mp8@802_g N_VDD_Mp8@802_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@801 N_OUT8_Mn8@801_d N_OUT7_Mn8@801_g N_VSS_Mn8@801_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@800 N_OUT8_Mn8@800_d N_OUT7_Mn8@800_g N_VSS_Mn8@800_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@801 N_OUT8_Mp8@801_d N_OUT7_Mp8@801_g N_VDD_Mp8@801_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@800 N_OUT8_Mp8@800_d N_OUT7_Mp8@800_g N_VDD_Mp8@800_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@799 N_OUT8_Mn8@799_d N_OUT7_Mn8@799_g N_VSS_Mn8@799_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@798 N_OUT8_Mn8@798_d N_OUT7_Mn8@798_g N_VSS_Mn8@798_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@799 N_OUT8_Mp8@799_d N_OUT7_Mp8@799_g N_VDD_Mp8@799_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@798 N_OUT8_Mp8@798_d N_OUT7_Mp8@798_g N_VDD_Mp8@798_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@797 N_OUT8_Mn8@797_d N_OUT7_Mn8@797_g N_VSS_Mn8@797_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@796 N_OUT8_Mn8@796_d N_OUT7_Mn8@796_g N_VSS_Mn8@796_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@797 N_OUT8_Mp8@797_d N_OUT7_Mp8@797_g N_VDD_Mp8@797_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@796 N_OUT8_Mp8@796_d N_OUT7_Mp8@796_g N_VDD_Mp8@796_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@795 N_OUT8_Mn8@795_d N_OUT7_Mn8@795_g N_VSS_Mn8@795_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@794 N_OUT8_Mn8@794_d N_OUT7_Mn8@794_g N_VSS_Mn8@794_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@795 N_OUT8_Mp8@795_d N_OUT7_Mp8@795_g N_VDD_Mp8@795_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@794 N_OUT8_Mp8@794_d N_OUT7_Mp8@794_g N_VDD_Mp8@794_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@793 N_OUT8_Mn8@793_d N_OUT7_Mn8@793_g N_VSS_Mn8@793_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@792 N_OUT8_Mn8@792_d N_OUT7_Mn8@792_g N_VSS_Mn8@792_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@793 N_OUT8_Mp8@793_d N_OUT7_Mp8@793_g N_VDD_Mp8@793_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@792 N_OUT8_Mp8@792_d N_OUT7_Mp8@792_g N_VDD_Mp8@792_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@791 N_OUT8_Mn8@791_d N_OUT7_Mn8@791_g N_VSS_Mn8@791_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@790 N_OUT8_Mn8@790_d N_OUT7_Mn8@790_g N_VSS_Mn8@790_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@791 N_OUT8_Mp8@791_d N_OUT7_Mp8@791_g N_VDD_Mp8@791_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@790 N_OUT8_Mp8@790_d N_OUT7_Mp8@790_g N_VDD_Mp8@790_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@789 N_OUT8_Mn8@789_d N_OUT7_Mn8@789_g N_VSS_Mn8@789_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@788 N_OUT8_Mn8@788_d N_OUT7_Mn8@788_g N_VSS_Mn8@788_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@789 N_OUT8_Mp8@789_d N_OUT7_Mp8@789_g N_VDD_Mp8@789_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@788 N_OUT8_Mp8@788_d N_OUT7_Mp8@788_g N_VDD_Mp8@788_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@787 N_OUT8_Mn8@787_d N_OUT7_Mn8@787_g N_VSS_Mn8@787_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@786 N_OUT8_Mn8@786_d N_OUT7_Mn8@786_g N_VSS_Mn8@786_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@787 N_OUT8_Mp8@787_d N_OUT7_Mp8@787_g N_VDD_Mp8@787_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@786 N_OUT8_Mp8@786_d N_OUT7_Mp8@786_g N_VDD_Mp8@786_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@785 N_OUT8_Mn8@785_d N_OUT7_Mn8@785_g N_VSS_Mn8@785_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@784 N_OUT8_Mn8@784_d N_OUT7_Mn8@784_g N_VSS_Mn8@784_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@785 N_OUT8_Mp8@785_d N_OUT7_Mp8@785_g N_VDD_Mp8@785_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@784 N_OUT8_Mp8@784_d N_OUT7_Mp8@784_g N_VDD_Mp8@784_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@783 N_OUT8_Mn8@783_d N_OUT7_Mn8@783_g N_VSS_Mn8@783_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@782 N_OUT8_Mn8@782_d N_OUT7_Mn8@782_g N_VSS_Mn8@782_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@783 N_OUT8_Mp8@783_d N_OUT7_Mp8@783_g N_VDD_Mp8@783_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@782 N_OUT8_Mp8@782_d N_OUT7_Mp8@782_g N_VDD_Mp8@782_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@781 N_OUT8_Mn8@781_d N_OUT7_Mn8@781_g N_VSS_Mn8@781_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@780 N_OUT8_Mn8@780_d N_OUT7_Mn8@780_g N_VSS_Mn8@780_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@781 N_OUT8_Mp8@781_d N_OUT7_Mp8@781_g N_VDD_Mp8@781_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@780 N_OUT8_Mp8@780_d N_OUT7_Mp8@780_g N_VDD_Mp8@780_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@779 N_OUT8_Mn8@779_d N_OUT7_Mn8@779_g N_VSS_Mn8@779_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@778 N_OUT8_Mn8@778_d N_OUT7_Mn8@778_g N_VSS_Mn8@778_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@779 N_OUT8_Mp8@779_d N_OUT7_Mp8@779_g N_VDD_Mp8@779_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@778 N_OUT8_Mp8@778_d N_OUT7_Mp8@778_g N_VDD_Mp8@778_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@777 N_OUT8_Mn8@777_d N_OUT7_Mn8@777_g N_VSS_Mn8@777_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@776 N_OUT8_Mn8@776_d N_OUT7_Mn8@776_g N_VSS_Mn8@776_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@777 N_OUT8_Mp8@777_d N_OUT7_Mp8@777_g N_VDD_Mp8@777_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@776 N_OUT8_Mp8@776_d N_OUT7_Mp8@776_g N_VDD_Mp8@776_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@775 N_OUT8_Mn8@775_d N_OUT7_Mn8@775_g N_VSS_Mn8@775_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@774 N_OUT8_Mn8@774_d N_OUT7_Mn8@774_g N_VSS_Mn8@774_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@775 N_OUT8_Mp8@775_d N_OUT7_Mp8@775_g N_VDD_Mp8@775_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@774 N_OUT8_Mp8@774_d N_OUT7_Mp8@774_g N_VDD_Mp8@774_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@773 N_OUT8_Mn8@773_d N_OUT7_Mn8@773_g N_VSS_Mn8@773_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@772 N_OUT8_Mn8@772_d N_OUT7_Mn8@772_g N_VSS_Mn8@772_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@773 N_OUT8_Mp8@773_d N_OUT7_Mp8@773_g N_VDD_Mp8@773_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@772 N_OUT8_Mp8@772_d N_OUT7_Mp8@772_g N_VDD_Mp8@772_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@771 N_OUT8_Mn8@771_d N_OUT7_Mn8@771_g N_VSS_Mn8@771_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@770 N_OUT8_Mn8@770_d N_OUT7_Mn8@770_g N_VSS_Mn8@770_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@771 N_OUT8_Mp8@771_d N_OUT7_Mp8@771_g N_VDD_Mp8@771_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@770 N_OUT8_Mp8@770_d N_OUT7_Mp8@770_g N_VDD_Mp8@770_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@769 N_OUT8_Mn8@769_d N_OUT7_Mn8@769_g N_VSS_Mn8@769_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@768 N_OUT8_Mn8@768_d N_OUT7_Mn8@768_g N_VSS_Mn8@768_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@769 N_OUT8_Mp8@769_d N_OUT7_Mp8@769_g N_VDD_Mp8@769_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@768 N_OUT8_Mp8@768_d N_OUT7_Mp8@768_g N_VDD_Mp8@768_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@767 N_OUT8_Mn8@767_d N_OUT7_Mn8@767_g N_VSS_Mn8@767_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@766 N_OUT8_Mn8@766_d N_OUT7_Mn8@766_g N_VSS_Mn8@766_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@767 N_OUT8_Mp8@767_d N_OUT7_Mp8@767_g N_VDD_Mp8@767_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@766 N_OUT8_Mp8@766_d N_OUT7_Mp8@766_g N_VDD_Mp8@766_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@765 N_OUT8_Mn8@765_d N_OUT7_Mn8@765_g N_VSS_Mn8@765_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@764 N_OUT8_Mn8@764_d N_OUT7_Mn8@764_g N_VSS_Mn8@764_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@765 N_OUT8_Mp8@765_d N_OUT7_Mp8@765_g N_VDD_Mp8@765_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@764 N_OUT8_Mp8@764_d N_OUT7_Mp8@764_g N_VDD_Mp8@764_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@763 N_OUT8_Mn8@763_d N_OUT7_Mn8@763_g N_VSS_Mn8@763_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@762 N_OUT8_Mn8@762_d N_OUT7_Mn8@762_g N_VSS_Mn8@762_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@763 N_OUT8_Mp8@763_d N_OUT7_Mp8@763_g N_VDD_Mp8@763_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@762 N_OUT8_Mp8@762_d N_OUT7_Mp8@762_g N_VDD_Mp8@762_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@761 N_OUT8_Mn8@761_d N_OUT7_Mn8@761_g N_VSS_Mn8@761_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@760 N_OUT8_Mn8@760_d N_OUT7_Mn8@760_g N_VSS_Mn8@760_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@761 N_OUT8_Mp8@761_d N_OUT7_Mp8@761_g N_VDD_Mp8@761_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@760 N_OUT8_Mp8@760_d N_OUT7_Mp8@760_g N_VDD_Mp8@760_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@759 N_OUT8_Mn8@759_d N_OUT7_Mn8@759_g N_VSS_Mn8@759_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@758 N_OUT8_Mn8@758_d N_OUT7_Mn8@758_g N_VSS_Mn8@758_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@759 N_OUT8_Mp8@759_d N_OUT7_Mp8@759_g N_VDD_Mp8@759_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@758 N_OUT8_Mp8@758_d N_OUT7_Mp8@758_g N_VDD_Mp8@758_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@757 N_OUT8_Mn8@757_d N_OUT7_Mn8@757_g N_VSS_Mn8@757_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@756 N_OUT8_Mn8@756_d N_OUT7_Mn8@756_g N_VSS_Mn8@756_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@757 N_OUT8_Mp8@757_d N_OUT7_Mp8@757_g N_VDD_Mp8@757_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@756 N_OUT8_Mp8@756_d N_OUT7_Mp8@756_g N_VDD_Mp8@756_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@755 N_OUT8_Mn8@755_d N_OUT7_Mn8@755_g N_VSS_Mn8@755_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@754 N_OUT8_Mn8@754_d N_OUT7_Mn8@754_g N_VSS_Mn8@754_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@755 N_OUT8_Mp8@755_d N_OUT7_Mp8@755_g N_VDD_Mp8@755_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@754 N_OUT8_Mp8@754_d N_OUT7_Mp8@754_g N_VDD_Mp8@754_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@753 N_OUT8_Mn8@753_d N_OUT7_Mn8@753_g N_VSS_Mn8@753_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@752 N_OUT8_Mn8@752_d N_OUT7_Mn8@752_g N_VSS_Mn8@752_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@753 N_OUT8_Mp8@753_d N_OUT7_Mp8@753_g N_VDD_Mp8@753_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@752 N_OUT8_Mp8@752_d N_OUT7_Mp8@752_g N_VDD_Mp8@752_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@751 N_OUT8_Mn8@751_d N_OUT7_Mn8@751_g N_VSS_Mn8@751_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@750 N_OUT8_Mn8@750_d N_OUT7_Mn8@750_g N_VSS_Mn8@750_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@751 N_OUT8_Mp8@751_d N_OUT7_Mp8@751_g N_VDD_Mp8@751_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@750 N_OUT8_Mp8@750_d N_OUT7_Mp8@750_g N_VDD_Mp8@750_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@749 N_OUT8_Mn8@749_d N_OUT7_Mn8@749_g N_VSS_Mn8@749_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@748 N_OUT8_Mn8@748_d N_OUT7_Mn8@748_g N_VSS_Mn8@748_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@749 N_OUT8_Mp8@749_d N_OUT7_Mp8@749_g N_VDD_Mp8@749_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@748 N_OUT8_Mp8@748_d N_OUT7_Mp8@748_g N_VDD_Mp8@748_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@747 N_OUT8_Mn8@747_d N_OUT7_Mn8@747_g N_VSS_Mn8@747_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@746 N_OUT8_Mn8@746_d N_OUT7_Mn8@746_g N_VSS_Mn8@746_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@747 N_OUT8_Mp8@747_d N_OUT7_Mp8@747_g N_VDD_Mp8@747_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@746 N_OUT8_Mp8@746_d N_OUT7_Mp8@746_g N_VDD_Mp8@746_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@745 N_OUT8_Mn8@745_d N_OUT7_Mn8@745_g N_VSS_Mn8@745_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@744 N_OUT8_Mn8@744_d N_OUT7_Mn8@744_g N_VSS_Mn8@744_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@745 N_OUT8_Mp8@745_d N_OUT7_Mp8@745_g N_VDD_Mp8@745_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@744 N_OUT8_Mp8@744_d N_OUT7_Mp8@744_g N_VDD_Mp8@744_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@743 N_OUT8_Mn8@743_d N_OUT7_Mn8@743_g N_VSS_Mn8@743_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@742 N_OUT8_Mn8@742_d N_OUT7_Mn8@742_g N_VSS_Mn8@742_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@743 N_OUT8_Mp8@743_d N_OUT7_Mp8@743_g N_VDD_Mp8@743_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@742 N_OUT8_Mp8@742_d N_OUT7_Mp8@742_g N_VDD_Mp8@742_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@741 N_OUT8_Mn8@741_d N_OUT7_Mn8@741_g N_VSS_Mn8@741_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@740 N_OUT8_Mn8@740_d N_OUT7_Mn8@740_g N_VSS_Mn8@740_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@741 N_OUT8_Mp8@741_d N_OUT7_Mp8@741_g N_VDD_Mp8@741_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@740 N_OUT8_Mp8@740_d N_OUT7_Mp8@740_g N_VDD_Mp8@740_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@739 N_OUT8_Mn8@739_d N_OUT7_Mn8@739_g N_VSS_Mn8@739_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@738 N_OUT8_Mn8@738_d N_OUT7_Mn8@738_g N_VSS_Mn8@738_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@739 N_OUT8_Mp8@739_d N_OUT7_Mp8@739_g N_VDD_Mp8@739_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@738 N_OUT8_Mp8@738_d N_OUT7_Mp8@738_g N_VDD_Mp8@738_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@737 N_OUT8_Mn8@737_d N_OUT7_Mn8@737_g N_VSS_Mn8@737_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@736 N_OUT8_Mn8@736_d N_OUT7_Mn8@736_g N_VSS_Mn8@736_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@737 N_OUT8_Mp8@737_d N_OUT7_Mp8@737_g N_VDD_Mp8@737_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@736 N_OUT8_Mp8@736_d N_OUT7_Mp8@736_g N_VDD_Mp8@736_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@735 N_OUT8_Mn8@735_d N_OUT7_Mn8@735_g N_VSS_Mn8@735_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@734 N_OUT8_Mn8@734_d N_OUT7_Mn8@734_g N_VSS_Mn8@734_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@735 N_OUT8_Mp8@735_d N_OUT7_Mp8@735_g N_VDD_Mp8@735_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@734 N_OUT8_Mp8@734_d N_OUT7_Mp8@734_g N_VDD_Mp8@734_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@733 N_OUT8_Mn8@733_d N_OUT7_Mn8@733_g N_VSS_Mn8@733_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@732 N_OUT8_Mn8@732_d N_OUT7_Mn8@732_g N_VSS_Mn8@732_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@733 N_OUT8_Mp8@733_d N_OUT7_Mp8@733_g N_VDD_Mp8@733_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@732 N_OUT8_Mp8@732_d N_OUT7_Mp8@732_g N_VDD_Mp8@732_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@731 N_OUT8_Mn8@731_d N_OUT7_Mn8@731_g N_VSS_Mn8@731_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@730 N_OUT8_Mn8@730_d N_OUT7_Mn8@730_g N_VSS_Mn8@730_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@731 N_OUT8_Mp8@731_d N_OUT7_Mp8@731_g N_VDD_Mp8@731_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@730 N_OUT8_Mp8@730_d N_OUT7_Mp8@730_g N_VDD_Mp8@730_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@729 N_OUT8_Mn8@729_d N_OUT7_Mn8@729_g N_VSS_Mn8@729_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@728 N_OUT8_Mn8@728_d N_OUT7_Mn8@728_g N_VSS_Mn8@728_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@729 N_OUT8_Mp8@729_d N_OUT7_Mp8@729_g N_VDD_Mp8@729_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@728 N_OUT8_Mp8@728_d N_OUT7_Mp8@728_g N_VDD_Mp8@728_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@727 N_OUT8_Mn8@727_d N_OUT7_Mn8@727_g N_VSS_Mn8@727_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@726 N_OUT8_Mn8@726_d N_OUT7_Mn8@726_g N_VSS_Mn8@726_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@727 N_OUT8_Mp8@727_d N_OUT7_Mp8@727_g N_VDD_Mp8@727_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@726 N_OUT8_Mp8@726_d N_OUT7_Mp8@726_g N_VDD_Mp8@726_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@725 N_OUT8_Mn8@725_d N_OUT7_Mn8@725_g N_VSS_Mn8@725_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@724 N_OUT8_Mn8@724_d N_OUT7_Mn8@724_g N_VSS_Mn8@724_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@725 N_OUT8_Mp8@725_d N_OUT7_Mp8@725_g N_VDD_Mp8@725_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@724 N_OUT8_Mp8@724_d N_OUT7_Mp8@724_g N_VDD_Mp8@724_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@723 N_OUT8_Mn8@723_d N_OUT7_Mn8@723_g N_VSS_Mn8@723_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@722 N_OUT8_Mn8@722_d N_OUT7_Mn8@722_g N_VSS_Mn8@722_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@723 N_OUT8_Mp8@723_d N_OUT7_Mp8@723_g N_VDD_Mp8@723_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@722 N_OUT8_Mp8@722_d N_OUT7_Mp8@722_g N_VDD_Mp8@722_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@721 N_OUT8_Mn8@721_d N_OUT7_Mn8@721_g N_VSS_Mn8@721_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@720 N_OUT8_Mn8@720_d N_OUT7_Mn8@720_g N_VSS_Mn8@720_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@721 N_OUT8_Mp8@721_d N_OUT7_Mp8@721_g N_VDD_Mp8@721_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@720 N_OUT8_Mp8@720_d N_OUT7_Mp8@720_g N_VDD_Mp8@720_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@719 N_OUT8_Mn8@719_d N_OUT7_Mn8@719_g N_VSS_Mn8@719_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@718 N_OUT8_Mn8@718_d N_OUT7_Mn8@718_g N_VSS_Mn8@718_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@719 N_OUT8_Mp8@719_d N_OUT7_Mp8@719_g N_VDD_Mp8@719_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@718 N_OUT8_Mp8@718_d N_OUT7_Mp8@718_g N_VDD_Mp8@718_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@717 N_OUT8_Mn8@717_d N_OUT7_Mn8@717_g N_VSS_Mn8@717_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@716 N_OUT8_Mn8@716_d N_OUT7_Mn8@716_g N_VSS_Mn8@716_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@717 N_OUT8_Mp8@717_d N_OUT7_Mp8@717_g N_VDD_Mp8@717_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@716 N_OUT8_Mp8@716_d N_OUT7_Mp8@716_g N_VDD_Mp8@716_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@715 N_OUT8_Mn8@715_d N_OUT7_Mn8@715_g N_VSS_Mn8@715_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@714 N_OUT8_Mn8@714_d N_OUT7_Mn8@714_g N_VSS_Mn8@714_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@715 N_OUT8_Mp8@715_d N_OUT7_Mp8@715_g N_VDD_Mp8@715_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@714 N_OUT8_Mp8@714_d N_OUT7_Mp8@714_g N_VDD_Mp8@714_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@713 N_OUT8_Mn8@713_d N_OUT7_Mn8@713_g N_VSS_Mn8@713_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@712 N_OUT8_Mn8@712_d N_OUT7_Mn8@712_g N_VSS_Mn8@712_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@713 N_OUT8_Mp8@713_d N_OUT7_Mp8@713_g N_VDD_Mp8@713_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@712 N_OUT8_Mp8@712_d N_OUT7_Mp8@712_g N_VDD_Mp8@712_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@711 N_OUT8_Mn8@711_d N_OUT7_Mn8@711_g N_VSS_Mn8@711_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@710 N_OUT8_Mn8@710_d N_OUT7_Mn8@710_g N_VSS_Mn8@710_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@711 N_OUT8_Mp8@711_d N_OUT7_Mp8@711_g N_VDD_Mp8@711_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@710 N_OUT8_Mp8@710_d N_OUT7_Mp8@710_g N_VDD_Mp8@710_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@709 N_OUT8_Mn8@709_d N_OUT7_Mn8@709_g N_VSS_Mn8@709_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@708 N_OUT8_Mn8@708_d N_OUT7_Mn8@708_g N_VSS_Mn8@708_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@709 N_OUT8_Mp8@709_d N_OUT7_Mp8@709_g N_VDD_Mp8@709_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@708 N_OUT8_Mp8@708_d N_OUT7_Mp8@708_g N_VDD_Mp8@708_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@707 N_OUT8_Mn8@707_d N_OUT7_Mn8@707_g N_VSS_Mn8@707_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@706 N_OUT8_Mn8@706_d N_OUT7_Mn8@706_g N_VSS_Mn8@706_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@707 N_OUT8_Mp8@707_d N_OUT7_Mp8@707_g N_VDD_Mp8@707_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@706 N_OUT8_Mp8@706_d N_OUT7_Mp8@706_g N_VDD_Mp8@706_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@705 N_OUT8_Mn8@705_d N_OUT7_Mn8@705_g N_VSS_Mn8@705_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@704 N_OUT8_Mn8@704_d N_OUT7_Mn8@704_g N_VSS_Mn8@704_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@705 N_OUT8_Mp8@705_d N_OUT7_Mp8@705_g N_VDD_Mp8@705_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@704 N_OUT8_Mp8@704_d N_OUT7_Mp8@704_g N_VDD_Mp8@704_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@703 N_OUT8_Mn8@703_d N_OUT7_Mn8@703_g N_VSS_Mn8@703_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@702 N_OUT8_Mn8@702_d N_OUT7_Mn8@702_g N_VSS_Mn8@702_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@703 N_OUT8_Mp8@703_d N_OUT7_Mp8@703_g N_VDD_Mp8@703_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@702 N_OUT8_Mp8@702_d N_OUT7_Mp8@702_g N_VDD_Mp8@702_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@701 N_OUT8_Mn8@701_d N_OUT7_Mn8@701_g N_VSS_Mn8@701_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@700 N_OUT8_Mn8@700_d N_OUT7_Mn8@700_g N_VSS_Mn8@700_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@701 N_OUT8_Mp8@701_d N_OUT7_Mp8@701_g N_VDD_Mp8@701_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@700 N_OUT8_Mp8@700_d N_OUT7_Mp8@700_g N_VDD_Mp8@700_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@699 N_OUT8_Mn8@699_d N_OUT7_Mn8@699_g N_VSS_Mn8@699_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@698 N_OUT8_Mn8@698_d N_OUT7_Mn8@698_g N_VSS_Mn8@698_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@699 N_OUT8_Mp8@699_d N_OUT7_Mp8@699_g N_VDD_Mp8@699_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@698 N_OUT8_Mp8@698_d N_OUT7_Mp8@698_g N_VDD_Mp8@698_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@697 N_OUT8_Mn8@697_d N_OUT7_Mn8@697_g N_VSS_Mn8@697_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@696 N_OUT8_Mn8@696_d N_OUT7_Mn8@696_g N_VSS_Mn8@696_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@697 N_OUT8_Mp8@697_d N_OUT7_Mp8@697_g N_VDD_Mp8@697_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@696 N_OUT8_Mp8@696_d N_OUT7_Mp8@696_g N_VDD_Mp8@696_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@695 N_OUT8_Mn8@695_d N_OUT7_Mn8@695_g N_VSS_Mn8@695_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@694 N_OUT8_Mn8@694_d N_OUT7_Mn8@694_g N_VSS_Mn8@694_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@695 N_OUT8_Mp8@695_d N_OUT7_Mp8@695_g N_VDD_Mp8@695_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@694 N_OUT8_Mp8@694_d N_OUT7_Mp8@694_g N_VDD_Mp8@694_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@693 N_OUT8_Mn8@693_d N_OUT7_Mn8@693_g N_VSS_Mn8@693_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@692 N_OUT8_Mn8@692_d N_OUT7_Mn8@692_g N_VSS_Mn8@692_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@693 N_OUT8_Mp8@693_d N_OUT7_Mp8@693_g N_VDD_Mp8@693_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@692 N_OUT8_Mp8@692_d N_OUT7_Mp8@692_g N_VDD_Mp8@692_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@691 N_OUT8_Mn8@691_d N_OUT7_Mn8@691_g N_VSS_Mn8@691_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@690 N_OUT8_Mn8@690_d N_OUT7_Mn8@690_g N_VSS_Mn8@690_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@691 N_OUT8_Mp8@691_d N_OUT7_Mp8@691_g N_VDD_Mp8@691_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@690 N_OUT8_Mp8@690_d N_OUT7_Mp8@690_g N_VDD_Mp8@690_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@689 N_OUT8_Mn8@689_d N_OUT7_Mn8@689_g N_VSS_Mn8@689_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@688 N_OUT8_Mn8@688_d N_OUT7_Mn8@688_g N_VSS_Mn8@688_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@689 N_OUT8_Mp8@689_d N_OUT7_Mp8@689_g N_VDD_Mp8@689_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@688 N_OUT8_Mp8@688_d N_OUT7_Mp8@688_g N_VDD_Mp8@688_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@687 N_OUT8_Mn8@687_d N_OUT7_Mn8@687_g N_VSS_Mn8@687_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@686 N_OUT8_Mn8@686_d N_OUT7_Mn8@686_g N_VSS_Mn8@686_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@687 N_OUT8_Mp8@687_d N_OUT7_Mp8@687_g N_VDD_Mp8@687_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@686 N_OUT8_Mp8@686_d N_OUT7_Mp8@686_g N_VDD_Mp8@686_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@685 N_OUT8_Mn8@685_d N_OUT7_Mn8@685_g N_VSS_Mn8@685_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@684 N_OUT8_Mn8@684_d N_OUT7_Mn8@684_g N_VSS_Mn8@684_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@685 N_OUT8_Mp8@685_d N_OUT7_Mp8@685_g N_VDD_Mp8@685_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@684 N_OUT8_Mp8@684_d N_OUT7_Mp8@684_g N_VDD_Mp8@684_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@683 N_OUT8_Mn8@683_d N_OUT7_Mn8@683_g N_VSS_Mn8@683_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@682 N_OUT8_Mn8@682_d N_OUT7_Mn8@682_g N_VSS_Mn8@682_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@683 N_OUT8_Mp8@683_d N_OUT7_Mp8@683_g N_VDD_Mp8@683_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@682 N_OUT8_Mp8@682_d N_OUT7_Mp8@682_g N_VDD_Mp8@682_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@681 N_OUT8_Mn8@681_d N_OUT7_Mn8@681_g N_VSS_Mn8@681_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@680 N_OUT8_Mn8@680_d N_OUT7_Mn8@680_g N_VSS_Mn8@680_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@681 N_OUT8_Mp8@681_d N_OUT7_Mp8@681_g N_VDD_Mp8@681_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@680 N_OUT8_Mp8@680_d N_OUT7_Mp8@680_g N_VDD_Mp8@680_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@679 N_OUT8_Mn8@679_d N_OUT7_Mn8@679_g N_VSS_Mn8@679_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@678 N_OUT8_Mn8@678_d N_OUT7_Mn8@678_g N_VSS_Mn8@678_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@679 N_OUT8_Mp8@679_d N_OUT7_Mp8@679_g N_VDD_Mp8@679_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@678 N_OUT8_Mp8@678_d N_OUT7_Mp8@678_g N_VDD_Mp8@678_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@677 N_OUT8_Mn8@677_d N_OUT7_Mn8@677_g N_VSS_Mn8@677_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@676 N_OUT8_Mn8@676_d N_OUT7_Mn8@676_g N_VSS_Mn8@676_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@677 N_OUT8_Mp8@677_d N_OUT7_Mp8@677_g N_VDD_Mp8@677_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@676 N_OUT8_Mp8@676_d N_OUT7_Mp8@676_g N_VDD_Mp8@676_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@675 N_OUT8_Mn8@675_d N_OUT7_Mn8@675_g N_VSS_Mn8@675_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@674 N_OUT8_Mn8@674_d N_OUT7_Mn8@674_g N_VSS_Mn8@674_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@675 N_OUT8_Mp8@675_d N_OUT7_Mp8@675_g N_VDD_Mp8@675_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@674 N_OUT8_Mp8@674_d N_OUT7_Mp8@674_g N_VDD_Mp8@674_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@673 N_OUT8_Mn8@673_d N_OUT7_Mn8@673_g N_VSS_Mn8@673_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@672 N_OUT8_Mn8@672_d N_OUT7_Mn8@672_g N_VSS_Mn8@672_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@673 N_OUT8_Mp8@673_d N_OUT7_Mp8@673_g N_VDD_Mp8@673_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@672 N_OUT8_Mp8@672_d N_OUT7_Mp8@672_g N_VDD_Mp8@672_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@671 N_OUT8_Mn8@671_d N_OUT7_Mn8@671_g N_VSS_Mn8@671_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@670 N_OUT8_Mn8@670_d N_OUT7_Mn8@670_g N_VSS_Mn8@670_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@671 N_OUT8_Mp8@671_d N_OUT7_Mp8@671_g N_VDD_Mp8@671_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@670 N_OUT8_Mp8@670_d N_OUT7_Mp8@670_g N_VDD_Mp8@670_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@669 N_OUT8_Mn8@669_d N_OUT7_Mn8@669_g N_VSS_Mn8@669_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@668 N_OUT8_Mn8@668_d N_OUT7_Mn8@668_g N_VSS_Mn8@668_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@669 N_OUT8_Mp8@669_d N_OUT7_Mp8@669_g N_VDD_Mp8@669_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@668 N_OUT8_Mp8@668_d N_OUT7_Mp8@668_g N_VDD_Mp8@668_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@667 N_OUT8_Mn8@667_d N_OUT7_Mn8@667_g N_VSS_Mn8@667_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@666 N_OUT8_Mn8@666_d N_OUT7_Mn8@666_g N_VSS_Mn8@666_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@667 N_OUT8_Mp8@667_d N_OUT7_Mp8@667_g N_VDD_Mp8@667_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@666 N_OUT8_Mp8@666_d N_OUT7_Mp8@666_g N_VDD_Mp8@666_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@665 N_OUT8_Mn8@665_d N_OUT7_Mn8@665_g N_VSS_Mn8@665_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@664 N_OUT8_Mn8@664_d N_OUT7_Mn8@664_g N_VSS_Mn8@664_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@665 N_OUT8_Mp8@665_d N_OUT7_Mp8@665_g N_VDD_Mp8@665_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@664 N_OUT8_Mp8@664_d N_OUT7_Mp8@664_g N_VDD_Mp8@664_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@663 N_OUT8_Mn8@663_d N_OUT7_Mn8@663_g N_VSS_Mn8@663_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@662 N_OUT8_Mn8@662_d N_OUT7_Mn8@662_g N_VSS_Mn8@662_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@663 N_OUT8_Mp8@663_d N_OUT7_Mp8@663_g N_VDD_Mp8@663_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@662 N_OUT8_Mp8@662_d N_OUT7_Mp8@662_g N_VDD_Mp8@662_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@661 N_OUT8_Mn8@661_d N_OUT7_Mn8@661_g N_VSS_Mn8@661_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@660 N_OUT8_Mn8@660_d N_OUT7_Mn8@660_g N_VSS_Mn8@660_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@661 N_OUT8_Mp8@661_d N_OUT7_Mp8@661_g N_VDD_Mp8@661_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@660 N_OUT8_Mp8@660_d N_OUT7_Mp8@660_g N_VDD_Mp8@660_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@659 N_OUT8_Mn8@659_d N_OUT7_Mn8@659_g N_VSS_Mn8@659_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@658 N_OUT8_Mn8@658_d N_OUT7_Mn8@658_g N_VSS_Mn8@658_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@659 N_OUT8_Mp8@659_d N_OUT7_Mp8@659_g N_VDD_Mp8@659_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@658 N_OUT8_Mp8@658_d N_OUT7_Mp8@658_g N_VDD_Mp8@658_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@657 N_OUT8_Mn8@657_d N_OUT7_Mn8@657_g N_VSS_Mn8@657_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@656 N_OUT8_Mn8@656_d N_OUT7_Mn8@656_g N_VSS_Mn8@656_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@657 N_OUT8_Mp8@657_d N_OUT7_Mp8@657_g N_VDD_Mp8@657_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@656 N_OUT8_Mp8@656_d N_OUT7_Mp8@656_g N_VDD_Mp8@656_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@655 N_OUT8_Mn8@655_d N_OUT7_Mn8@655_g N_VSS_Mn8@655_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@654 N_OUT8_Mn8@654_d N_OUT7_Mn8@654_g N_VSS_Mn8@654_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@655 N_OUT8_Mp8@655_d N_OUT7_Mp8@655_g N_VDD_Mp8@655_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@654 N_OUT8_Mp8@654_d N_OUT7_Mp8@654_g N_VDD_Mp8@654_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@653 N_OUT8_Mn8@653_d N_OUT7_Mn8@653_g N_VSS_Mn8@653_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@652 N_OUT8_Mn8@652_d N_OUT7_Mn8@652_g N_VSS_Mn8@652_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@653 N_OUT8_Mp8@653_d N_OUT7_Mp8@653_g N_VDD_Mp8@653_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@652 N_OUT8_Mp8@652_d N_OUT7_Mp8@652_g N_VDD_Mp8@652_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@651 N_OUT8_Mn8@651_d N_OUT7_Mn8@651_g N_VSS_Mn8@651_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@650 N_OUT8_Mn8@650_d N_OUT7_Mn8@650_g N_VSS_Mn8@650_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@651 N_OUT8_Mp8@651_d N_OUT7_Mp8@651_g N_VDD_Mp8@651_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@650 N_OUT8_Mp8@650_d N_OUT7_Mp8@650_g N_VDD_Mp8@650_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@649 N_OUT8_Mn8@649_d N_OUT7_Mn8@649_g N_VSS_Mn8@649_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@648 N_OUT8_Mn8@648_d N_OUT7_Mn8@648_g N_VSS_Mn8@648_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@649 N_OUT8_Mp8@649_d N_OUT7_Mp8@649_g N_VDD_Mp8@649_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@648 N_OUT8_Mp8@648_d N_OUT7_Mp8@648_g N_VDD_Mp8@648_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@647 N_OUT8_Mn8@647_d N_OUT7_Mn8@647_g N_VSS_Mn8@647_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@646 N_OUT8_Mn8@646_d N_OUT7_Mn8@646_g N_VSS_Mn8@646_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@647 N_OUT8_Mp8@647_d N_OUT7_Mp8@647_g N_VDD_Mp8@647_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@646 N_OUT8_Mp8@646_d N_OUT7_Mp8@646_g N_VDD_Mp8@646_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@645 N_OUT8_Mn8@645_d N_OUT7_Mn8@645_g N_VSS_Mn8@645_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@644 N_OUT8_Mn8@644_d N_OUT7_Mn8@644_g N_VSS_Mn8@644_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@645 N_OUT8_Mp8@645_d N_OUT7_Mp8@645_g N_VDD_Mp8@645_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@644 N_OUT8_Mp8@644_d N_OUT7_Mp8@644_g N_VDD_Mp8@644_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@643 N_OUT8_Mn8@643_d N_OUT7_Mn8@643_g N_VSS_Mn8@643_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@642 N_OUT8_Mn8@642_d N_OUT7_Mn8@642_g N_VSS_Mn8@642_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@643 N_OUT8_Mp8@643_d N_OUT7_Mp8@643_g N_VDD_Mp8@643_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@642 N_OUT8_Mp8@642_d N_OUT7_Mp8@642_g N_VDD_Mp8@642_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@641 N_OUT8_Mn8@641_d N_OUT7_Mn8@641_g N_VSS_Mn8@641_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@640 N_OUT8_Mn8@640_d N_OUT7_Mn8@640_g N_VSS_Mn8@640_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@641 N_OUT8_Mp8@641_d N_OUT7_Mp8@641_g N_VDD_Mp8@641_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@640 N_OUT8_Mp8@640_d N_OUT7_Mp8@640_g N_VDD_Mp8@640_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@639 N_OUT8_Mn8@639_d N_OUT7_Mn8@639_g N_VSS_Mn8@639_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@638 N_OUT8_Mn8@638_d N_OUT7_Mn8@638_g N_VSS_Mn8@638_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@639 N_OUT8_Mp8@639_d N_OUT7_Mp8@639_g N_VDD_Mp8@639_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@638 N_OUT8_Mp8@638_d N_OUT7_Mp8@638_g N_VDD_Mp8@638_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@637 N_OUT8_Mn8@637_d N_OUT7_Mn8@637_g N_VSS_Mn8@637_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@636 N_OUT8_Mn8@636_d N_OUT7_Mn8@636_g N_VSS_Mn8@636_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@637 N_OUT8_Mp8@637_d N_OUT7_Mp8@637_g N_VDD_Mp8@637_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@636 N_OUT8_Mp8@636_d N_OUT7_Mp8@636_g N_VDD_Mp8@636_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@635 N_OUT8_Mn8@635_d N_OUT7_Mn8@635_g N_VSS_Mn8@635_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@634 N_OUT8_Mn8@634_d N_OUT7_Mn8@634_g N_VSS_Mn8@634_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@635 N_OUT8_Mp8@635_d N_OUT7_Mp8@635_g N_VDD_Mp8@635_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@634 N_OUT8_Mp8@634_d N_OUT7_Mp8@634_g N_VDD_Mp8@634_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@633 N_OUT8_Mn8@633_d N_OUT7_Mn8@633_g N_VSS_Mn8@633_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@632 N_OUT8_Mn8@632_d N_OUT7_Mn8@632_g N_VSS_Mn8@632_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@633 N_OUT8_Mp8@633_d N_OUT7_Mp8@633_g N_VDD_Mp8@633_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@632 N_OUT8_Mp8@632_d N_OUT7_Mp8@632_g N_VDD_Mp8@632_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@631 N_OUT8_Mn8@631_d N_OUT7_Mn8@631_g N_VSS_Mn8@631_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@630 N_OUT8_Mn8@630_d N_OUT7_Mn8@630_g N_VSS_Mn8@630_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@631 N_OUT8_Mp8@631_d N_OUT7_Mp8@631_g N_VDD_Mp8@631_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@630 N_OUT8_Mp8@630_d N_OUT7_Mp8@630_g N_VDD_Mp8@630_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@629 N_OUT8_Mn8@629_d N_OUT7_Mn8@629_g N_VSS_Mn8@629_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@628 N_OUT8_Mn8@628_d N_OUT7_Mn8@628_g N_VSS_Mn8@628_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@629 N_OUT8_Mp8@629_d N_OUT7_Mp8@629_g N_VDD_Mp8@629_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@628 N_OUT8_Mp8@628_d N_OUT7_Mp8@628_g N_VDD_Mp8@628_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@627 N_OUT8_Mn8@627_d N_OUT7_Mn8@627_g N_VSS_Mn8@627_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@626 N_OUT8_Mn8@626_d N_OUT7_Mn8@626_g N_VSS_Mn8@626_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@627 N_OUT8_Mp8@627_d N_OUT7_Mp8@627_g N_VDD_Mp8@627_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@626 N_OUT8_Mp8@626_d N_OUT7_Mp8@626_g N_VDD_Mp8@626_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@625 N_OUT8_Mn8@625_d N_OUT7_Mn8@625_g N_VSS_Mn8@625_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@624 N_OUT8_Mn8@624_d N_OUT7_Mn8@624_g N_VSS_Mn8@624_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@625 N_OUT8_Mp8@625_d N_OUT7_Mp8@625_g N_VDD_Mp8@625_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@624 N_OUT8_Mp8@624_d N_OUT7_Mp8@624_g N_VDD_Mp8@624_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@623 N_OUT8_Mn8@623_d N_OUT7_Mn8@623_g N_VSS_Mn8@623_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@622 N_OUT8_Mn8@622_d N_OUT7_Mn8@622_g N_VSS_Mn8@622_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@623 N_OUT8_Mp8@623_d N_OUT7_Mp8@623_g N_VDD_Mp8@623_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@622 N_OUT8_Mp8@622_d N_OUT7_Mp8@622_g N_VDD_Mp8@622_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@621 N_OUT8_Mn8@621_d N_OUT7_Mn8@621_g N_VSS_Mn8@621_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@620 N_OUT8_Mn8@620_d N_OUT7_Mn8@620_g N_VSS_Mn8@620_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@621 N_OUT8_Mp8@621_d N_OUT7_Mp8@621_g N_VDD_Mp8@621_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@620 N_OUT8_Mp8@620_d N_OUT7_Mp8@620_g N_VDD_Mp8@620_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@619 N_OUT8_Mn8@619_d N_OUT7_Mn8@619_g N_VSS_Mn8@619_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@618 N_OUT8_Mn8@618_d N_OUT7_Mn8@618_g N_VSS_Mn8@618_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@619 N_OUT8_Mp8@619_d N_OUT7_Mp8@619_g N_VDD_Mp8@619_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@618 N_OUT8_Mp8@618_d N_OUT7_Mp8@618_g N_VDD_Mp8@618_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@617 N_OUT8_Mn8@617_d N_OUT7_Mn8@617_g N_VSS_Mn8@617_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@616 N_OUT8_Mn8@616_d N_OUT7_Mn8@616_g N_VSS_Mn8@616_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@617 N_OUT8_Mp8@617_d N_OUT7_Mp8@617_g N_VDD_Mp8@617_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@616 N_OUT8_Mp8@616_d N_OUT7_Mp8@616_g N_VDD_Mp8@616_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@615 N_OUT8_Mn8@615_d N_OUT7_Mn8@615_g N_VSS_Mn8@615_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@614 N_OUT8_Mn8@614_d N_OUT7_Mn8@614_g N_VSS_Mn8@614_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@615 N_OUT8_Mp8@615_d N_OUT7_Mp8@615_g N_VDD_Mp8@615_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@614 N_OUT8_Mp8@614_d N_OUT7_Mp8@614_g N_VDD_Mp8@614_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@613 N_OUT8_Mn8@613_d N_OUT7_Mn8@613_g N_VSS_Mn8@613_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@612 N_OUT8_Mn8@612_d N_OUT7_Mn8@612_g N_VSS_Mn8@612_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@613 N_OUT8_Mp8@613_d N_OUT7_Mp8@613_g N_VDD_Mp8@613_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@612 N_OUT8_Mp8@612_d N_OUT7_Mp8@612_g N_VDD_Mp8@612_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@611 N_OUT8_Mn8@611_d N_OUT7_Mn8@611_g N_VSS_Mn8@611_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@610 N_OUT8_Mn8@610_d N_OUT7_Mn8@610_g N_VSS_Mn8@610_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@611 N_OUT8_Mp8@611_d N_OUT7_Mp8@611_g N_VDD_Mp8@611_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@610 N_OUT8_Mp8@610_d N_OUT7_Mp8@610_g N_VDD_Mp8@610_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@609 N_OUT8_Mn8@609_d N_OUT7_Mn8@609_g N_VSS_Mn8@609_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@608 N_OUT8_Mn8@608_d N_OUT7_Mn8@608_g N_VSS_Mn8@608_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@609 N_OUT8_Mp8@609_d N_OUT7_Mp8@609_g N_VDD_Mp8@609_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@608 N_OUT8_Mp8@608_d N_OUT7_Mp8@608_g N_VDD_Mp8@608_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@607 N_OUT8_Mn8@607_d N_OUT7_Mn8@607_g N_VSS_Mn8@607_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@606 N_OUT8_Mn8@606_d N_OUT7_Mn8@606_g N_VSS_Mn8@606_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@607 N_OUT8_Mp8@607_d N_OUT7_Mp8@607_g N_VDD_Mp8@607_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@606 N_OUT8_Mp8@606_d N_OUT7_Mp8@606_g N_VDD_Mp8@606_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@605 N_OUT8_Mn8@605_d N_OUT7_Mn8@605_g N_VSS_Mn8@605_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@604 N_OUT8_Mn8@604_d N_OUT7_Mn8@604_g N_VSS_Mn8@604_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@605 N_OUT8_Mp8@605_d N_OUT7_Mp8@605_g N_VDD_Mp8@605_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@604 N_OUT8_Mp8@604_d N_OUT7_Mp8@604_g N_VDD_Mp8@604_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@603 N_OUT8_Mn8@603_d N_OUT7_Mn8@603_g N_VSS_Mn8@603_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@602 N_OUT8_Mn8@602_d N_OUT7_Mn8@602_g N_VSS_Mn8@602_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@603 N_OUT8_Mp8@603_d N_OUT7_Mp8@603_g N_VDD_Mp8@603_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@602 N_OUT8_Mp8@602_d N_OUT7_Mp8@602_g N_VDD_Mp8@602_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@601 N_OUT8_Mn8@601_d N_OUT7_Mn8@601_g N_VSS_Mn8@601_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@600 N_OUT8_Mn8@600_d N_OUT7_Mn8@600_g N_VSS_Mn8@600_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@601 N_OUT8_Mp8@601_d N_OUT7_Mp8@601_g N_VDD_Mp8@601_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@600 N_OUT8_Mp8@600_d N_OUT7_Mp8@600_g N_VDD_Mp8@600_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@599 N_OUT8_Mn8@599_d N_OUT7_Mn8@599_g N_VSS_Mn8@599_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@598 N_OUT8_Mn8@598_d N_OUT7_Mn8@598_g N_VSS_Mn8@598_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@599 N_OUT8_Mp8@599_d N_OUT7_Mp8@599_g N_VDD_Mp8@599_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@598 N_OUT8_Mp8@598_d N_OUT7_Mp8@598_g N_VDD_Mp8@598_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@597 N_OUT8_Mn8@597_d N_OUT7_Mn8@597_g N_VSS_Mn8@597_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@596 N_OUT8_Mn8@596_d N_OUT7_Mn8@596_g N_VSS_Mn8@596_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@597 N_OUT8_Mp8@597_d N_OUT7_Mp8@597_g N_VDD_Mp8@597_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@596 N_OUT8_Mp8@596_d N_OUT7_Mp8@596_g N_VDD_Mp8@596_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@595 N_OUT8_Mn8@595_d N_OUT7_Mn8@595_g N_VSS_Mn8@595_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@594 N_OUT8_Mn8@594_d N_OUT7_Mn8@594_g N_VSS_Mn8@594_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@595 N_OUT8_Mp8@595_d N_OUT7_Mp8@595_g N_VDD_Mp8@595_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@594 N_OUT8_Mp8@594_d N_OUT7_Mp8@594_g N_VDD_Mp8@594_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@593 N_OUT8_Mn8@593_d N_OUT7_Mn8@593_g N_VSS_Mn8@593_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@592 N_OUT8_Mn8@592_d N_OUT7_Mn8@592_g N_VSS_Mn8@592_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@593 N_OUT8_Mp8@593_d N_OUT7_Mp8@593_g N_VDD_Mp8@593_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@592 N_OUT8_Mp8@592_d N_OUT7_Mp8@592_g N_VDD_Mp8@592_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@591 N_OUT8_Mn8@591_d N_OUT7_Mn8@591_g N_VSS_Mn8@591_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@590 N_OUT8_Mn8@590_d N_OUT7_Mn8@590_g N_VSS_Mn8@590_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@591 N_OUT8_Mp8@591_d N_OUT7_Mp8@591_g N_VDD_Mp8@591_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@590 N_OUT8_Mp8@590_d N_OUT7_Mp8@590_g N_VDD_Mp8@590_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@589 N_OUT8_Mn8@589_d N_OUT7_Mn8@589_g N_VSS_Mn8@589_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@588 N_OUT8_Mn8@588_d N_OUT7_Mn8@588_g N_VSS_Mn8@588_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@589 N_OUT8_Mp8@589_d N_OUT7_Mp8@589_g N_VDD_Mp8@589_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@588 N_OUT8_Mp8@588_d N_OUT7_Mp8@588_g N_VDD_Mp8@588_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@587 N_OUT8_Mn8@587_d N_OUT7_Mn8@587_g N_VSS_Mn8@587_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@586 N_OUT8_Mn8@586_d N_OUT7_Mn8@586_g N_VSS_Mn8@586_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@587 N_OUT8_Mp8@587_d N_OUT7_Mp8@587_g N_VDD_Mp8@587_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@586 N_OUT8_Mp8@586_d N_OUT7_Mp8@586_g N_VDD_Mp8@586_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@585 N_OUT8_Mn8@585_d N_OUT7_Mn8@585_g N_VSS_Mn8@585_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@584 N_OUT8_Mn8@584_d N_OUT7_Mn8@584_g N_VSS_Mn8@584_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@585 N_OUT8_Mp8@585_d N_OUT7_Mp8@585_g N_VDD_Mp8@585_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@584 N_OUT8_Mp8@584_d N_OUT7_Mp8@584_g N_VDD_Mp8@584_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@583 N_OUT8_Mn8@583_d N_OUT7_Mn8@583_g N_VSS_Mn8@583_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@582 N_OUT8_Mn8@582_d N_OUT7_Mn8@582_g N_VSS_Mn8@582_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@583 N_OUT8_Mp8@583_d N_OUT7_Mp8@583_g N_VDD_Mp8@583_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@582 N_OUT8_Mp8@582_d N_OUT7_Mp8@582_g N_VDD_Mp8@582_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@581 N_OUT8_Mn8@581_d N_OUT7_Mn8@581_g N_VSS_Mn8@581_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@580 N_OUT8_Mn8@580_d N_OUT7_Mn8@580_g N_VSS_Mn8@580_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@581 N_OUT8_Mp8@581_d N_OUT7_Mp8@581_g N_VDD_Mp8@581_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@580 N_OUT8_Mp8@580_d N_OUT7_Mp8@580_g N_VDD_Mp8@580_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@579 N_OUT8_Mn8@579_d N_OUT7_Mn8@579_g N_VSS_Mn8@579_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@578 N_OUT8_Mn8@578_d N_OUT7_Mn8@578_g N_VSS_Mn8@578_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@579 N_OUT8_Mp8@579_d N_OUT7_Mp8@579_g N_VDD_Mp8@579_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@578 N_OUT8_Mp8@578_d N_OUT7_Mp8@578_g N_VDD_Mp8@578_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@577 N_OUT8_Mn8@577_d N_OUT7_Mn8@577_g N_VSS_Mn8@577_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@576 N_OUT8_Mn8@576_d N_OUT7_Mn8@576_g N_VSS_Mn8@576_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@577 N_OUT8_Mp8@577_d N_OUT7_Mp8@577_g N_VDD_Mp8@577_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@576 N_OUT8_Mp8@576_d N_OUT7_Mp8@576_g N_VDD_Mp8@576_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@575 N_OUT8_Mn8@575_d N_OUT7_Mn8@575_g N_VSS_Mn8@575_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@574 N_OUT8_Mn8@574_d N_OUT7_Mn8@574_g N_VSS_Mn8@574_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@575 N_OUT8_Mp8@575_d N_OUT7_Mp8@575_g N_VDD_Mp8@575_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@574 N_OUT8_Mp8@574_d N_OUT7_Mp8@574_g N_VDD_Mp8@574_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@573 N_OUT8_Mn8@573_d N_OUT7_Mn8@573_g N_VSS_Mn8@573_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@572 N_OUT8_Mn8@572_d N_OUT7_Mn8@572_g N_VSS_Mn8@572_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@573 N_OUT8_Mp8@573_d N_OUT7_Mp8@573_g N_VDD_Mp8@573_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@572 N_OUT8_Mp8@572_d N_OUT7_Mp8@572_g N_VDD_Mp8@572_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@571 N_OUT8_Mn8@571_d N_OUT7_Mn8@571_g N_VSS_Mn8@571_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@570 N_OUT8_Mn8@570_d N_OUT7_Mn8@570_g N_VSS_Mn8@570_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@571 N_OUT8_Mp8@571_d N_OUT7_Mp8@571_g N_VDD_Mp8@571_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@570 N_OUT8_Mp8@570_d N_OUT7_Mp8@570_g N_VDD_Mp8@570_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@569 N_OUT8_Mn8@569_d N_OUT7_Mn8@569_g N_VSS_Mn8@569_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@568 N_OUT8_Mn8@568_d N_OUT7_Mn8@568_g N_VSS_Mn8@568_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@569 N_OUT8_Mp8@569_d N_OUT7_Mp8@569_g N_VDD_Mp8@569_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@568 N_OUT8_Mp8@568_d N_OUT7_Mp8@568_g N_VDD_Mp8@568_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@567 N_OUT8_Mn8@567_d N_OUT7_Mn8@567_g N_VSS_Mn8@567_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@566 N_OUT8_Mn8@566_d N_OUT7_Mn8@566_g N_VSS_Mn8@566_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@567 N_OUT8_Mp8@567_d N_OUT7_Mp8@567_g N_VDD_Mp8@567_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@566 N_OUT8_Mp8@566_d N_OUT7_Mp8@566_g N_VDD_Mp8@566_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@565 N_OUT8_Mn8@565_d N_OUT7_Mn8@565_g N_VSS_Mn8@565_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@564 N_OUT8_Mn8@564_d N_OUT7_Mn8@564_g N_VSS_Mn8@564_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@565 N_OUT8_Mp8@565_d N_OUT7_Mp8@565_g N_VDD_Mp8@565_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@564 N_OUT8_Mp8@564_d N_OUT7_Mp8@564_g N_VDD_Mp8@564_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@563 N_OUT8_Mn8@563_d N_OUT7_Mn8@563_g N_VSS_Mn8@563_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@562 N_OUT8_Mn8@562_d N_OUT7_Mn8@562_g N_VSS_Mn8@562_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@563 N_OUT8_Mp8@563_d N_OUT7_Mp8@563_g N_VDD_Mp8@563_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@562 N_OUT8_Mp8@562_d N_OUT7_Mp8@562_g N_VDD_Mp8@562_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@561 N_OUT8_Mn8@561_d N_OUT7_Mn8@561_g N_VSS_Mn8@561_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@560 N_OUT8_Mn8@560_d N_OUT7_Mn8@560_g N_VSS_Mn8@560_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@561 N_OUT8_Mp8@561_d N_OUT7_Mp8@561_g N_VDD_Mp8@561_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@560 N_OUT8_Mp8@560_d N_OUT7_Mp8@560_g N_VDD_Mp8@560_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@559 N_OUT8_Mn8@559_d N_OUT7_Mn8@559_g N_VSS_Mn8@559_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@558 N_OUT8_Mn8@558_d N_OUT7_Mn8@558_g N_VSS_Mn8@558_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@559 N_OUT8_Mp8@559_d N_OUT7_Mp8@559_g N_VDD_Mp8@559_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@558 N_OUT8_Mp8@558_d N_OUT7_Mp8@558_g N_VDD_Mp8@558_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@557 N_OUT8_Mn8@557_d N_OUT7_Mn8@557_g N_VSS_Mn8@557_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@556 N_OUT8_Mn8@556_d N_OUT7_Mn8@556_g N_VSS_Mn8@556_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@557 N_OUT8_Mp8@557_d N_OUT7_Mp8@557_g N_VDD_Mp8@557_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@556 N_OUT8_Mp8@556_d N_OUT7_Mp8@556_g N_VDD_Mp8@556_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@555 N_OUT8_Mn8@555_d N_OUT7_Mn8@555_g N_VSS_Mn8@555_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@554 N_OUT8_Mn8@554_d N_OUT7_Mn8@554_g N_VSS_Mn8@554_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@555 N_OUT8_Mp8@555_d N_OUT7_Mp8@555_g N_VDD_Mp8@555_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@554 N_OUT8_Mp8@554_d N_OUT7_Mp8@554_g N_VDD_Mp8@554_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@553 N_OUT8_Mn8@553_d N_OUT7_Mn8@553_g N_VSS_Mn8@553_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@552 N_OUT8_Mn8@552_d N_OUT7_Mn8@552_g N_VSS_Mn8@552_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@553 N_OUT8_Mp8@553_d N_OUT7_Mp8@553_g N_VDD_Mp8@553_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@552 N_OUT8_Mp8@552_d N_OUT7_Mp8@552_g N_VDD_Mp8@552_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@551 N_OUT8_Mn8@551_d N_OUT7_Mn8@551_g N_VSS_Mn8@551_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@550 N_OUT8_Mn8@550_d N_OUT7_Mn8@550_g N_VSS_Mn8@550_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@551 N_OUT8_Mp8@551_d N_OUT7_Mp8@551_g N_VDD_Mp8@551_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@550 N_OUT8_Mp8@550_d N_OUT7_Mp8@550_g N_VDD_Mp8@550_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@549 N_OUT8_Mn8@549_d N_OUT7_Mn8@549_g N_VSS_Mn8@549_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@548 N_OUT8_Mn8@548_d N_OUT7_Mn8@548_g N_VSS_Mn8@548_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@549 N_OUT8_Mp8@549_d N_OUT7_Mp8@549_g N_VDD_Mp8@549_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@548 N_OUT8_Mp8@548_d N_OUT7_Mp8@548_g N_VDD_Mp8@548_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@547 N_OUT8_Mn8@547_d N_OUT7_Mn8@547_g N_VSS_Mn8@547_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@546 N_OUT8_Mn8@546_d N_OUT7_Mn8@546_g N_VSS_Mn8@546_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@547 N_OUT8_Mp8@547_d N_OUT7_Mp8@547_g N_VDD_Mp8@547_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@546 N_OUT8_Mp8@546_d N_OUT7_Mp8@546_g N_VDD_Mp8@546_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@545 N_OUT8_Mn8@545_d N_OUT7_Mn8@545_g N_VSS_Mn8@545_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@544 N_OUT8_Mn8@544_d N_OUT7_Mn8@544_g N_VSS_Mn8@544_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@545 N_OUT8_Mp8@545_d N_OUT7_Mp8@545_g N_VDD_Mp8@545_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@544 N_OUT8_Mp8@544_d N_OUT7_Mp8@544_g N_VDD_Mp8@544_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@543 N_OUT8_Mn8@543_d N_OUT7_Mn8@543_g N_VSS_Mn8@543_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@542 N_OUT8_Mn8@542_d N_OUT7_Mn8@542_g N_VSS_Mn8@542_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@543 N_OUT8_Mp8@543_d N_OUT7_Mp8@543_g N_VDD_Mp8@543_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@542 N_OUT8_Mp8@542_d N_OUT7_Mp8@542_g N_VDD_Mp8@542_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@541 N_OUT8_Mn8@541_d N_OUT7_Mn8@541_g N_VSS_Mn8@541_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@540 N_OUT8_Mn8@540_d N_OUT7_Mn8@540_g N_VSS_Mn8@540_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@541 N_OUT8_Mp8@541_d N_OUT7_Mp8@541_g N_VDD_Mp8@541_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@540 N_OUT8_Mp8@540_d N_OUT7_Mp8@540_g N_VDD_Mp8@540_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@539 N_OUT8_Mn8@539_d N_OUT7_Mn8@539_g N_VSS_Mn8@539_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@538 N_OUT8_Mn8@538_d N_OUT7_Mn8@538_g N_VSS_Mn8@538_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@539 N_OUT8_Mp8@539_d N_OUT7_Mp8@539_g N_VDD_Mp8@539_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@538 N_OUT8_Mp8@538_d N_OUT7_Mp8@538_g N_VDD_Mp8@538_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@537 N_OUT8_Mn8@537_d N_OUT7_Mn8@537_g N_VSS_Mn8@537_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@536 N_OUT8_Mn8@536_d N_OUT7_Mn8@536_g N_VSS_Mn8@536_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@537 N_OUT8_Mp8@537_d N_OUT7_Mp8@537_g N_VDD_Mp8@537_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@536 N_OUT8_Mp8@536_d N_OUT7_Mp8@536_g N_VDD_Mp8@536_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@535 N_OUT8_Mn8@535_d N_OUT7_Mn8@535_g N_VSS_Mn8@535_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@534 N_OUT8_Mn8@534_d N_OUT7_Mn8@534_g N_VSS_Mn8@534_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@535 N_OUT8_Mp8@535_d N_OUT7_Mp8@535_g N_VDD_Mp8@535_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@534 N_OUT8_Mp8@534_d N_OUT7_Mp8@534_g N_VDD_Mp8@534_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@533 N_OUT8_Mn8@533_d N_OUT7_Mn8@533_g N_VSS_Mn8@533_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@532 N_OUT8_Mn8@532_d N_OUT7_Mn8@532_g N_VSS_Mn8@532_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@533 N_OUT8_Mp8@533_d N_OUT7_Mp8@533_g N_VDD_Mp8@533_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@532 N_OUT8_Mp8@532_d N_OUT7_Mp8@532_g N_VDD_Mp8@532_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@531 N_OUT8_Mn8@531_d N_OUT7_Mn8@531_g N_VSS_Mn8@531_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@530 N_OUT8_Mn8@530_d N_OUT7_Mn8@530_g N_VSS_Mn8@530_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@531 N_OUT8_Mp8@531_d N_OUT7_Mp8@531_g N_VDD_Mp8@531_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@530 N_OUT8_Mp8@530_d N_OUT7_Mp8@530_g N_VDD_Mp8@530_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@529 N_OUT8_Mn8@529_d N_OUT7_Mn8@529_g N_VSS_Mn8@529_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@528 N_OUT8_Mn8@528_d N_OUT7_Mn8@528_g N_VSS_Mn8@528_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@529 N_OUT8_Mp8@529_d N_OUT7_Mp8@529_g N_VDD_Mp8@529_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@528 N_OUT8_Mp8@528_d N_OUT7_Mp8@528_g N_VDD_Mp8@528_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@527 N_OUT8_Mn8@527_d N_OUT7_Mn8@527_g N_VSS_Mn8@527_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@526 N_OUT8_Mn8@526_d N_OUT7_Mn8@526_g N_VSS_Mn8@526_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@527 N_OUT8_Mp8@527_d N_OUT7_Mp8@527_g N_VDD_Mp8@527_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@526 N_OUT8_Mp8@526_d N_OUT7_Mp8@526_g N_VDD_Mp8@526_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@525 N_OUT8_Mn8@525_d N_OUT7_Mn8@525_g N_VSS_Mn8@525_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@524 N_OUT8_Mn8@524_d N_OUT7_Mn8@524_g N_VSS_Mn8@524_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@525 N_OUT8_Mp8@525_d N_OUT7_Mp8@525_g N_VDD_Mp8@525_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@524 N_OUT8_Mp8@524_d N_OUT7_Mp8@524_g N_VDD_Mp8@524_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@523 N_OUT8_Mn8@523_d N_OUT7_Mn8@523_g N_VSS_Mn8@523_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@522 N_OUT8_Mn8@522_d N_OUT7_Mn8@522_g N_VSS_Mn8@522_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@523 N_OUT8_Mp8@523_d N_OUT7_Mp8@523_g N_VDD_Mp8@523_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@522 N_OUT8_Mp8@522_d N_OUT7_Mp8@522_g N_VDD_Mp8@522_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@521 N_OUT8_Mn8@521_d N_OUT7_Mn8@521_g N_VSS_Mn8@521_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@520 N_OUT8_Mn8@520_d N_OUT7_Mn8@520_g N_VSS_Mn8@520_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@521 N_OUT8_Mp8@521_d N_OUT7_Mp8@521_g N_VDD_Mp8@521_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@520 N_OUT8_Mp8@520_d N_OUT7_Mp8@520_g N_VDD_Mp8@520_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@519 N_OUT8_Mn8@519_d N_OUT7_Mn8@519_g N_VSS_Mn8@519_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@518 N_OUT8_Mn8@518_d N_OUT7_Mn8@518_g N_VSS_Mn8@518_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@519 N_OUT8_Mp8@519_d N_OUT7_Mp8@519_g N_VDD_Mp8@519_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@518 N_OUT8_Mp8@518_d N_OUT7_Mp8@518_g N_VDD_Mp8@518_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@517 N_OUT8_Mn8@517_d N_OUT7_Mn8@517_g N_VSS_Mn8@517_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@516 N_OUT8_Mn8@516_d N_OUT7_Mn8@516_g N_VSS_Mn8@516_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@517 N_OUT8_Mp8@517_d N_OUT7_Mp8@517_g N_VDD_Mp8@517_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@516 N_OUT8_Mp8@516_d N_OUT7_Mp8@516_g N_VDD_Mp8@516_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@515 N_OUT8_Mn8@515_d N_OUT7_Mn8@515_g N_VSS_Mn8@515_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@514 N_OUT8_Mn8@514_d N_OUT7_Mn8@514_g N_VSS_Mn8@514_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@515 N_OUT8_Mp8@515_d N_OUT7_Mp8@515_g N_VDD_Mp8@515_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@514 N_OUT8_Mp8@514_d N_OUT7_Mp8@514_g N_VDD_Mp8@514_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@513 N_OUT8_Mn8@513_d N_OUT7_Mn8@513_g N_VSS_Mn8@513_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@512 N_OUT8_Mn8@512_d N_OUT7_Mn8@512_g N_VSS_Mn8@512_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@513 N_OUT8_Mp8@513_d N_OUT7_Mp8@513_g N_VDD_Mp8@513_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@512 N_OUT8_Mp8@512_d N_OUT7_Mp8@512_g N_VDD_Mp8@512_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@511 N_OUT8_Mn8@511_d N_OUT7_Mn8@511_g N_VSS_Mn8@511_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@510 N_OUT8_Mn8@510_d N_OUT7_Mn8@510_g N_VSS_Mn8@510_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@511 N_OUT8_Mp8@511_d N_OUT7_Mp8@511_g N_VDD_Mp8@511_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@510 N_OUT8_Mp8@510_d N_OUT7_Mp8@510_g N_VDD_Mp8@510_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@509 N_OUT8_Mn8@509_d N_OUT7_Mn8@509_g N_VSS_Mn8@509_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@508 N_OUT8_Mn8@508_d N_OUT7_Mn8@508_g N_VSS_Mn8@508_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@509 N_OUT8_Mp8@509_d N_OUT7_Mp8@509_g N_VDD_Mp8@509_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@508 N_OUT8_Mp8@508_d N_OUT7_Mp8@508_g N_VDD_Mp8@508_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@507 N_OUT8_Mn8@507_d N_OUT7_Mn8@507_g N_VSS_Mn8@507_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@506 N_OUT8_Mn8@506_d N_OUT7_Mn8@506_g N_VSS_Mn8@506_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@507 N_OUT8_Mp8@507_d N_OUT7_Mp8@507_g N_VDD_Mp8@507_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@506 N_OUT8_Mp8@506_d N_OUT7_Mp8@506_g N_VDD_Mp8@506_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@505 N_OUT8_Mn8@505_d N_OUT7_Mn8@505_g N_VSS_Mn8@505_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@504 N_OUT8_Mn8@504_d N_OUT7_Mn8@504_g N_VSS_Mn8@504_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@505 N_OUT8_Mp8@505_d N_OUT7_Mp8@505_g N_VDD_Mp8@505_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@504 N_OUT8_Mp8@504_d N_OUT7_Mp8@504_g N_VDD_Mp8@504_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@503 N_OUT8_Mn8@503_d N_OUT7_Mn8@503_g N_VSS_Mn8@503_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@502 N_OUT8_Mn8@502_d N_OUT7_Mn8@502_g N_VSS_Mn8@502_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@503 N_OUT8_Mp8@503_d N_OUT7_Mp8@503_g N_VDD_Mp8@503_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@502 N_OUT8_Mp8@502_d N_OUT7_Mp8@502_g N_VDD_Mp8@502_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@501 N_OUT8_Mn8@501_d N_OUT7_Mn8@501_g N_VSS_Mn8@501_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@500 N_OUT8_Mn8@500_d N_OUT7_Mn8@500_g N_VSS_Mn8@500_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@501 N_OUT8_Mp8@501_d N_OUT7_Mp8@501_g N_VDD_Mp8@501_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@500 N_OUT8_Mp8@500_d N_OUT7_Mp8@500_g N_VDD_Mp8@500_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@499 N_OUT8_Mn8@499_d N_OUT7_Mn8@499_g N_VSS_Mn8@499_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@498 N_OUT8_Mn8@498_d N_OUT7_Mn8@498_g N_VSS_Mn8@498_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@499 N_OUT8_Mp8@499_d N_OUT7_Mp8@499_g N_VDD_Mp8@499_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@498 N_OUT8_Mp8@498_d N_OUT7_Mp8@498_g N_VDD_Mp8@498_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@497 N_OUT8_Mn8@497_d N_OUT7_Mn8@497_g N_VSS_Mn8@497_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@496 N_OUT8_Mn8@496_d N_OUT7_Mn8@496_g N_VSS_Mn8@496_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@497 N_OUT8_Mp8@497_d N_OUT7_Mp8@497_g N_VDD_Mp8@497_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@496 N_OUT8_Mp8@496_d N_OUT7_Mp8@496_g N_VDD_Mp8@496_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@495 N_OUT8_Mn8@495_d N_OUT7_Mn8@495_g N_VSS_Mn8@495_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@494 N_OUT8_Mn8@494_d N_OUT7_Mn8@494_g N_VSS_Mn8@494_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@495 N_OUT8_Mp8@495_d N_OUT7_Mp8@495_g N_VDD_Mp8@495_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@494 N_OUT8_Mp8@494_d N_OUT7_Mp8@494_g N_VDD_Mp8@494_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@493 N_OUT8_Mn8@493_d N_OUT7_Mn8@493_g N_VSS_Mn8@493_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@492 N_OUT8_Mn8@492_d N_OUT7_Mn8@492_g N_VSS_Mn8@492_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@493 N_OUT8_Mp8@493_d N_OUT7_Mp8@493_g N_VDD_Mp8@493_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@492 N_OUT8_Mp8@492_d N_OUT7_Mp8@492_g N_VDD_Mp8@492_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@491 N_OUT8_Mn8@491_d N_OUT7_Mn8@491_g N_VSS_Mn8@491_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@490 N_OUT8_Mn8@490_d N_OUT7_Mn8@490_g N_VSS_Mn8@490_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@491 N_OUT8_Mp8@491_d N_OUT7_Mp8@491_g N_VDD_Mp8@491_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@490 N_OUT8_Mp8@490_d N_OUT7_Mp8@490_g N_VDD_Mp8@490_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@489 N_OUT8_Mn8@489_d N_OUT7_Mn8@489_g N_VSS_Mn8@489_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@488 N_OUT8_Mn8@488_d N_OUT7_Mn8@488_g N_VSS_Mn8@488_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@489 N_OUT8_Mp8@489_d N_OUT7_Mp8@489_g N_VDD_Mp8@489_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@488 N_OUT8_Mp8@488_d N_OUT7_Mp8@488_g N_VDD_Mp8@488_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@487 N_OUT8_Mn8@487_d N_OUT7_Mn8@487_g N_VSS_Mn8@487_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@486 N_OUT8_Mn8@486_d N_OUT7_Mn8@486_g N_VSS_Mn8@486_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@487 N_OUT8_Mp8@487_d N_OUT7_Mp8@487_g N_VDD_Mp8@487_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@486 N_OUT8_Mp8@486_d N_OUT7_Mp8@486_g N_VDD_Mp8@486_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@485 N_OUT8_Mn8@485_d N_OUT7_Mn8@485_g N_VSS_Mn8@485_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@484 N_OUT8_Mn8@484_d N_OUT7_Mn8@484_g N_VSS_Mn8@484_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@485 N_OUT8_Mp8@485_d N_OUT7_Mp8@485_g N_VDD_Mp8@485_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@484 N_OUT8_Mp8@484_d N_OUT7_Mp8@484_g N_VDD_Mp8@484_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@483 N_OUT8_Mn8@483_d N_OUT7_Mn8@483_g N_VSS_Mn8@483_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@482 N_OUT8_Mn8@482_d N_OUT7_Mn8@482_g N_VSS_Mn8@482_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@483 N_OUT8_Mp8@483_d N_OUT7_Mp8@483_g N_VDD_Mp8@483_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@482 N_OUT8_Mp8@482_d N_OUT7_Mp8@482_g N_VDD_Mp8@482_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@481 N_OUT8_Mn8@481_d N_OUT7_Mn8@481_g N_VSS_Mn8@481_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@480 N_OUT8_Mn8@480_d N_OUT7_Mn8@480_g N_VSS_Mn8@480_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@481 N_OUT8_Mp8@481_d N_OUT7_Mp8@481_g N_VDD_Mp8@481_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@480 N_OUT8_Mp8@480_d N_OUT7_Mp8@480_g N_VDD_Mp8@480_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@479 N_OUT8_Mn8@479_d N_OUT7_Mn8@479_g N_VSS_Mn8@479_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@478 N_OUT8_Mn8@478_d N_OUT7_Mn8@478_g N_VSS_Mn8@478_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@479 N_OUT8_Mp8@479_d N_OUT7_Mp8@479_g N_VDD_Mp8@479_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@478 N_OUT8_Mp8@478_d N_OUT7_Mp8@478_g N_VDD_Mp8@478_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@477 N_OUT8_Mn8@477_d N_OUT7_Mn8@477_g N_VSS_Mn8@477_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@476 N_OUT8_Mn8@476_d N_OUT7_Mn8@476_g N_VSS_Mn8@476_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@477 N_OUT8_Mp8@477_d N_OUT7_Mp8@477_g N_VDD_Mp8@477_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@476 N_OUT8_Mp8@476_d N_OUT7_Mp8@476_g N_VDD_Mp8@476_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@475 N_OUT8_Mn8@475_d N_OUT7_Mn8@475_g N_VSS_Mn8@475_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@474 N_OUT8_Mn8@474_d N_OUT7_Mn8@474_g N_VSS_Mn8@474_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@475 N_OUT8_Mp8@475_d N_OUT7_Mp8@475_g N_VDD_Mp8@475_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@474 N_OUT8_Mp8@474_d N_OUT7_Mp8@474_g N_VDD_Mp8@474_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@473 N_OUT8_Mn8@473_d N_OUT7_Mn8@473_g N_VSS_Mn8@473_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@472 N_OUT8_Mn8@472_d N_OUT7_Mn8@472_g N_VSS_Mn8@472_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@473 N_OUT8_Mp8@473_d N_OUT7_Mp8@473_g N_VDD_Mp8@473_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@472 N_OUT8_Mp8@472_d N_OUT7_Mp8@472_g N_VDD_Mp8@472_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@471 N_OUT8_Mn8@471_d N_OUT7_Mn8@471_g N_VSS_Mn8@471_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@470 N_OUT8_Mn8@470_d N_OUT7_Mn8@470_g N_VSS_Mn8@470_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@471 N_OUT8_Mp8@471_d N_OUT7_Mp8@471_g N_VDD_Mp8@471_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@470 N_OUT8_Mp8@470_d N_OUT7_Mp8@470_g N_VDD_Mp8@470_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@469 N_OUT8_Mn8@469_d N_OUT7_Mn8@469_g N_VSS_Mn8@469_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@468 N_OUT8_Mn8@468_d N_OUT7_Mn8@468_g N_VSS_Mn8@468_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@469 N_OUT8_Mp8@469_d N_OUT7_Mp8@469_g N_VDD_Mp8@469_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@468 N_OUT8_Mp8@468_d N_OUT7_Mp8@468_g N_VDD_Mp8@468_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@467 N_OUT8_Mn8@467_d N_OUT7_Mn8@467_g N_VSS_Mn8@467_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@466 N_OUT8_Mn8@466_d N_OUT7_Mn8@466_g N_VSS_Mn8@466_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@467 N_OUT8_Mp8@467_d N_OUT7_Mp8@467_g N_VDD_Mp8@467_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@466 N_OUT8_Mp8@466_d N_OUT7_Mp8@466_g N_VDD_Mp8@466_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@465 N_OUT8_Mn8@465_d N_OUT7_Mn8@465_g N_VSS_Mn8@465_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@464 N_OUT8_Mn8@464_d N_OUT7_Mn8@464_g N_VSS_Mn8@464_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@465 N_OUT8_Mp8@465_d N_OUT7_Mp8@465_g N_VDD_Mp8@465_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@464 N_OUT8_Mp8@464_d N_OUT7_Mp8@464_g N_VDD_Mp8@464_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@463 N_OUT8_Mn8@463_d N_OUT7_Mn8@463_g N_VSS_Mn8@463_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@462 N_OUT8_Mn8@462_d N_OUT7_Mn8@462_g N_VSS_Mn8@462_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@463 N_OUT8_Mp8@463_d N_OUT7_Mp8@463_g N_VDD_Mp8@463_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@462 N_OUT8_Mp8@462_d N_OUT7_Mp8@462_g N_VDD_Mp8@462_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@461 N_OUT8_Mn8@461_d N_OUT7_Mn8@461_g N_VSS_Mn8@461_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@460 N_OUT8_Mn8@460_d N_OUT7_Mn8@460_g N_VSS_Mn8@460_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@461 N_OUT8_Mp8@461_d N_OUT7_Mp8@461_g N_VDD_Mp8@461_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@460 N_OUT8_Mp8@460_d N_OUT7_Mp8@460_g N_VDD_Mp8@460_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@459 N_OUT8_Mn8@459_d N_OUT7_Mn8@459_g N_VSS_Mn8@459_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@458 N_OUT8_Mn8@458_d N_OUT7_Mn8@458_g N_VSS_Mn8@458_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@459 N_OUT8_Mp8@459_d N_OUT7_Mp8@459_g N_VDD_Mp8@459_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@458 N_OUT8_Mp8@458_d N_OUT7_Mp8@458_g N_VDD_Mp8@458_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@457 N_OUT8_Mn8@457_d N_OUT7_Mn8@457_g N_VSS_Mn8@457_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@456 N_OUT8_Mn8@456_d N_OUT7_Mn8@456_g N_VSS_Mn8@456_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@457 N_OUT8_Mp8@457_d N_OUT7_Mp8@457_g N_VDD_Mp8@457_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@456 N_OUT8_Mp8@456_d N_OUT7_Mp8@456_g N_VDD_Mp8@456_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@455 N_OUT8_Mn8@455_d N_OUT7_Mn8@455_g N_VSS_Mn8@455_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@454 N_OUT8_Mn8@454_d N_OUT7_Mn8@454_g N_VSS_Mn8@454_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@455 N_OUT8_Mp8@455_d N_OUT7_Mp8@455_g N_VDD_Mp8@455_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@454 N_OUT8_Mp8@454_d N_OUT7_Mp8@454_g N_VDD_Mp8@454_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@453 N_OUT8_Mn8@453_d N_OUT7_Mn8@453_g N_VSS_Mn8@453_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@452 N_OUT8_Mn8@452_d N_OUT7_Mn8@452_g N_VSS_Mn8@452_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@453 N_OUT8_Mp8@453_d N_OUT7_Mp8@453_g N_VDD_Mp8@453_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@452 N_OUT8_Mp8@452_d N_OUT7_Mp8@452_g N_VDD_Mp8@452_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@451 N_OUT8_Mn8@451_d N_OUT7_Mn8@451_g N_VSS_Mn8@451_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@450 N_OUT8_Mn8@450_d N_OUT7_Mn8@450_g N_VSS_Mn8@450_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@451 N_OUT8_Mp8@451_d N_OUT7_Mp8@451_g N_VDD_Mp8@451_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@450 N_OUT8_Mp8@450_d N_OUT7_Mp8@450_g N_VDD_Mp8@450_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@449 N_OUT8_Mn8@449_d N_OUT7_Mn8@449_g N_VSS_Mn8@449_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@448 N_OUT8_Mn8@448_d N_OUT7_Mn8@448_g N_VSS_Mn8@448_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@449 N_OUT8_Mp8@449_d N_OUT7_Mp8@449_g N_VDD_Mp8@449_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@448 N_OUT8_Mp8@448_d N_OUT7_Mp8@448_g N_VDD_Mp8@448_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@447 N_OUT8_Mn8@447_d N_OUT7_Mn8@447_g N_VSS_Mn8@447_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@446 N_OUT8_Mn8@446_d N_OUT7_Mn8@446_g N_VSS_Mn8@446_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@447 N_OUT8_Mp8@447_d N_OUT7_Mp8@447_g N_VDD_Mp8@447_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@446 N_OUT8_Mp8@446_d N_OUT7_Mp8@446_g N_VDD_Mp8@446_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@445 N_OUT8_Mn8@445_d N_OUT7_Mn8@445_g N_VSS_Mn8@445_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@444 N_OUT8_Mn8@444_d N_OUT7_Mn8@444_g N_VSS_Mn8@444_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@445 N_OUT8_Mp8@445_d N_OUT7_Mp8@445_g N_VDD_Mp8@445_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@444 N_OUT8_Mp8@444_d N_OUT7_Mp8@444_g N_VDD_Mp8@444_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@443 N_OUT8_Mn8@443_d N_OUT7_Mn8@443_g N_VSS_Mn8@443_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@442 N_OUT8_Mn8@442_d N_OUT7_Mn8@442_g N_VSS_Mn8@442_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@443 N_OUT8_Mp8@443_d N_OUT7_Mp8@443_g N_VDD_Mp8@443_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@442 N_OUT8_Mp8@442_d N_OUT7_Mp8@442_g N_VDD_Mp8@442_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@441 N_OUT8_Mn8@441_d N_OUT7_Mn8@441_g N_VSS_Mn8@441_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@440 N_OUT8_Mn8@440_d N_OUT7_Mn8@440_g N_VSS_Mn8@440_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@441 N_OUT8_Mp8@441_d N_OUT7_Mp8@441_g N_VDD_Mp8@441_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@440 N_OUT8_Mp8@440_d N_OUT7_Mp8@440_g N_VDD_Mp8@440_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@439 N_OUT8_Mn8@439_d N_OUT7_Mn8@439_g N_VSS_Mn8@439_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@438 N_OUT8_Mn8@438_d N_OUT7_Mn8@438_g N_VSS_Mn8@438_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@439 N_OUT8_Mp8@439_d N_OUT7_Mp8@439_g N_VDD_Mp8@439_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@438 N_OUT8_Mp8@438_d N_OUT7_Mp8@438_g N_VDD_Mp8@438_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@437 N_OUT8_Mn8@437_d N_OUT7_Mn8@437_g N_VSS_Mn8@437_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@436 N_OUT8_Mn8@436_d N_OUT7_Mn8@436_g N_VSS_Mn8@436_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@437 N_OUT8_Mp8@437_d N_OUT7_Mp8@437_g N_VDD_Mp8@437_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@436 N_OUT8_Mp8@436_d N_OUT7_Mp8@436_g N_VDD_Mp8@436_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@435 N_OUT8_Mn8@435_d N_OUT7_Mn8@435_g N_VSS_Mn8@435_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@434 N_OUT8_Mn8@434_d N_OUT7_Mn8@434_g N_VSS_Mn8@434_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@435 N_OUT8_Mp8@435_d N_OUT7_Mp8@435_g N_VDD_Mp8@435_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@434 N_OUT8_Mp8@434_d N_OUT7_Mp8@434_g N_VDD_Mp8@434_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@433 N_OUT8_Mn8@433_d N_OUT7_Mn8@433_g N_VSS_Mn8@433_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@432 N_OUT8_Mn8@432_d N_OUT7_Mn8@432_g N_VSS_Mn8@432_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@433 N_OUT8_Mp8@433_d N_OUT7_Mp8@433_g N_VDD_Mp8@433_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@432 N_OUT8_Mp8@432_d N_OUT7_Mp8@432_g N_VDD_Mp8@432_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@431 N_OUT8_Mn8@431_d N_OUT7_Mn8@431_g N_VSS_Mn8@431_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@430 N_OUT8_Mn8@430_d N_OUT7_Mn8@430_g N_VSS_Mn8@430_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@431 N_OUT8_Mp8@431_d N_OUT7_Mp8@431_g N_VDD_Mp8@431_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@430 N_OUT8_Mp8@430_d N_OUT7_Mp8@430_g N_VDD_Mp8@430_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@429 N_OUT8_Mn8@429_d N_OUT7_Mn8@429_g N_VSS_Mn8@429_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@428 N_OUT8_Mn8@428_d N_OUT7_Mn8@428_g N_VSS_Mn8@428_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@429 N_OUT8_Mp8@429_d N_OUT7_Mp8@429_g N_VDD_Mp8@429_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@428 N_OUT8_Mp8@428_d N_OUT7_Mp8@428_g N_VDD_Mp8@428_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@427 N_OUT8_Mn8@427_d N_OUT7_Mn8@427_g N_VSS_Mn8@427_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@426 N_OUT8_Mn8@426_d N_OUT7_Mn8@426_g N_VSS_Mn8@426_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@427 N_OUT8_Mp8@427_d N_OUT7_Mp8@427_g N_VDD_Mp8@427_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@426 N_OUT8_Mp8@426_d N_OUT7_Mp8@426_g N_VDD_Mp8@426_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@425 N_OUT8_Mn8@425_d N_OUT7_Mn8@425_g N_VSS_Mn8@425_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@424 N_OUT8_Mn8@424_d N_OUT7_Mn8@424_g N_VSS_Mn8@424_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@425 N_OUT8_Mp8@425_d N_OUT7_Mp8@425_g N_VDD_Mp8@425_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@424 N_OUT8_Mp8@424_d N_OUT7_Mp8@424_g N_VDD_Mp8@424_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@423 N_OUT8_Mn8@423_d N_OUT7_Mn8@423_g N_VSS_Mn8@423_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@422 N_OUT8_Mn8@422_d N_OUT7_Mn8@422_g N_VSS_Mn8@422_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@423 N_OUT8_Mp8@423_d N_OUT7_Mp8@423_g N_VDD_Mp8@423_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@422 N_OUT8_Mp8@422_d N_OUT7_Mp8@422_g N_VDD_Mp8@422_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@421 N_OUT8_Mn8@421_d N_OUT7_Mn8@421_g N_VSS_Mn8@421_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@420 N_OUT8_Mn8@420_d N_OUT7_Mn8@420_g N_VSS_Mn8@420_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@421 N_OUT8_Mp8@421_d N_OUT7_Mp8@421_g N_VDD_Mp8@421_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@420 N_OUT8_Mp8@420_d N_OUT7_Mp8@420_g N_VDD_Mp8@420_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@419 N_OUT8_Mn8@419_d N_OUT7_Mn8@419_g N_VSS_Mn8@419_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@418 N_OUT8_Mn8@418_d N_OUT7_Mn8@418_g N_VSS_Mn8@418_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@419 N_OUT8_Mp8@419_d N_OUT7_Mp8@419_g N_VDD_Mp8@419_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@418 N_OUT8_Mp8@418_d N_OUT7_Mp8@418_g N_VDD_Mp8@418_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@417 N_OUT8_Mn8@417_d N_OUT7_Mn8@417_g N_VSS_Mn8@417_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@416 N_OUT8_Mn8@416_d N_OUT7_Mn8@416_g N_VSS_Mn8@416_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@417 N_OUT8_Mp8@417_d N_OUT7_Mp8@417_g N_VDD_Mp8@417_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@416 N_OUT8_Mp8@416_d N_OUT7_Mp8@416_g N_VDD_Mp8@416_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@415 N_OUT8_Mn8@415_d N_OUT7_Mn8@415_g N_VSS_Mn8@415_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@414 N_OUT8_Mn8@414_d N_OUT7_Mn8@414_g N_VSS_Mn8@414_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@415 N_OUT8_Mp8@415_d N_OUT7_Mp8@415_g N_VDD_Mp8@415_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@414 N_OUT8_Mp8@414_d N_OUT7_Mp8@414_g N_VDD_Mp8@414_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@413 N_OUT8_Mn8@413_d N_OUT7_Mn8@413_g N_VSS_Mn8@413_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@412 N_OUT8_Mn8@412_d N_OUT7_Mn8@412_g N_VSS_Mn8@412_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@413 N_OUT8_Mp8@413_d N_OUT7_Mp8@413_g N_VDD_Mp8@413_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@412 N_OUT8_Mp8@412_d N_OUT7_Mp8@412_g N_VDD_Mp8@412_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@411 N_OUT8_Mn8@411_d N_OUT7_Mn8@411_g N_VSS_Mn8@411_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@410 N_OUT8_Mn8@410_d N_OUT7_Mn8@410_g N_VSS_Mn8@410_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@411 N_OUT8_Mp8@411_d N_OUT7_Mp8@411_g N_VDD_Mp8@411_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@410 N_OUT8_Mp8@410_d N_OUT7_Mp8@410_g N_VDD_Mp8@410_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@409 N_OUT8_Mn8@409_d N_OUT7_Mn8@409_g N_VSS_Mn8@409_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@408 N_OUT8_Mn8@408_d N_OUT7_Mn8@408_g N_VSS_Mn8@408_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@409 N_OUT8_Mp8@409_d N_OUT7_Mp8@409_g N_VDD_Mp8@409_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@408 N_OUT8_Mp8@408_d N_OUT7_Mp8@408_g N_VDD_Mp8@408_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@407 N_OUT8_Mn8@407_d N_OUT7_Mn8@407_g N_VSS_Mn8@407_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@406 N_OUT8_Mn8@406_d N_OUT7_Mn8@406_g N_VSS_Mn8@406_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@407 N_OUT8_Mp8@407_d N_OUT7_Mp8@407_g N_VDD_Mp8@407_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@406 N_OUT8_Mp8@406_d N_OUT7_Mp8@406_g N_VDD_Mp8@406_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@405 N_OUT8_Mn8@405_d N_OUT7_Mn8@405_g N_VSS_Mn8@405_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@404 N_OUT8_Mn8@404_d N_OUT7_Mn8@404_g N_VSS_Mn8@404_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@405 N_OUT8_Mp8@405_d N_OUT7_Mp8@405_g N_VDD_Mp8@405_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@404 N_OUT8_Mp8@404_d N_OUT7_Mp8@404_g N_VDD_Mp8@404_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@403 N_OUT8_Mn8@403_d N_OUT7_Mn8@403_g N_VSS_Mn8@403_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@402 N_OUT8_Mn8@402_d N_OUT7_Mn8@402_g N_VSS_Mn8@402_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@403 N_OUT8_Mp8@403_d N_OUT7_Mp8@403_g N_VDD_Mp8@403_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@402 N_OUT8_Mp8@402_d N_OUT7_Mp8@402_g N_VDD_Mp8@402_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@401 N_OUT8_Mn8@401_d N_OUT7_Mn8@401_g N_VSS_Mn8@401_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@400 N_OUT8_Mn8@400_d N_OUT7_Mn8@400_g N_VSS_Mn8@400_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@401 N_OUT8_Mp8@401_d N_OUT7_Mp8@401_g N_VDD_Mp8@401_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@400 N_OUT8_Mp8@400_d N_OUT7_Mp8@400_g N_VDD_Mp8@400_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@399 N_OUT8_Mn8@399_d N_OUT7_Mn8@399_g N_VSS_Mn8@399_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@398 N_OUT8_Mn8@398_d N_OUT7_Mn8@398_g N_VSS_Mn8@398_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@399 N_OUT8_Mp8@399_d N_OUT7_Mp8@399_g N_VDD_Mp8@399_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@398 N_OUT8_Mp8@398_d N_OUT7_Mp8@398_g N_VDD_Mp8@398_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@397 N_OUT8_Mn8@397_d N_OUT7_Mn8@397_g N_VSS_Mn8@397_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@396 N_OUT8_Mn8@396_d N_OUT7_Mn8@396_g N_VSS_Mn8@396_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@397 N_OUT8_Mp8@397_d N_OUT7_Mp8@397_g N_VDD_Mp8@397_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@396 N_OUT8_Mp8@396_d N_OUT7_Mp8@396_g N_VDD_Mp8@396_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@395 N_OUT8_Mn8@395_d N_OUT7_Mn8@395_g N_VSS_Mn8@395_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@394 N_OUT8_Mn8@394_d N_OUT7_Mn8@394_g N_VSS_Mn8@394_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@395 N_OUT8_Mp8@395_d N_OUT7_Mp8@395_g N_VDD_Mp8@395_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@394 N_OUT8_Mp8@394_d N_OUT7_Mp8@394_g N_VDD_Mp8@394_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@393 N_OUT8_Mn8@393_d N_OUT7_Mn8@393_g N_VSS_Mn8@393_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@392 N_OUT8_Mn8@392_d N_OUT7_Mn8@392_g N_VSS_Mn8@392_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@393 N_OUT8_Mp8@393_d N_OUT7_Mp8@393_g N_VDD_Mp8@393_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@392 N_OUT8_Mp8@392_d N_OUT7_Mp8@392_g N_VDD_Mp8@392_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@391 N_OUT8_Mn8@391_d N_OUT7_Mn8@391_g N_VSS_Mn8@391_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@390 N_OUT8_Mn8@390_d N_OUT7_Mn8@390_g N_VSS_Mn8@390_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@391 N_OUT8_Mp8@391_d N_OUT7_Mp8@391_g N_VDD_Mp8@391_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@390 N_OUT8_Mp8@390_d N_OUT7_Mp8@390_g N_VDD_Mp8@390_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@389 N_OUT8_Mn8@389_d N_OUT7_Mn8@389_g N_VSS_Mn8@389_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@388 N_OUT8_Mn8@388_d N_OUT7_Mn8@388_g N_VSS_Mn8@388_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@389 N_OUT8_Mp8@389_d N_OUT7_Mp8@389_g N_VDD_Mp8@389_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@388 N_OUT8_Mp8@388_d N_OUT7_Mp8@388_g N_VDD_Mp8@388_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@387 N_OUT8_Mn8@387_d N_OUT7_Mn8@387_g N_VSS_Mn8@387_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@386 N_OUT8_Mn8@386_d N_OUT7_Mn8@386_g N_VSS_Mn8@386_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@387 N_OUT8_Mp8@387_d N_OUT7_Mp8@387_g N_VDD_Mp8@387_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@386 N_OUT8_Mp8@386_d N_OUT7_Mp8@386_g N_VDD_Mp8@386_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@385 N_OUT8_Mn8@385_d N_OUT7_Mn8@385_g N_VSS_Mn8@385_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@384 N_OUT8_Mn8@384_d N_OUT7_Mn8@384_g N_VSS_Mn8@384_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@385 N_OUT8_Mp8@385_d N_OUT7_Mp8@385_g N_VDD_Mp8@385_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@384 N_OUT8_Mp8@384_d N_OUT7_Mp8@384_g N_VDD_Mp8@384_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@383 N_OUT8_Mn8@383_d N_OUT7_Mn8@383_g N_VSS_Mn8@383_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@382 N_OUT8_Mn8@382_d N_OUT7_Mn8@382_g N_VSS_Mn8@382_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@383 N_OUT8_Mp8@383_d N_OUT7_Mp8@383_g N_VDD_Mp8@383_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@382 N_OUT8_Mp8@382_d N_OUT7_Mp8@382_g N_VDD_Mp8@382_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@381 N_OUT8_Mn8@381_d N_OUT7_Mn8@381_g N_VSS_Mn8@381_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@380 N_OUT8_Mn8@380_d N_OUT7_Mn8@380_g N_VSS_Mn8@380_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@381 N_OUT8_Mp8@381_d N_OUT7_Mp8@381_g N_VDD_Mp8@381_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@380 N_OUT8_Mp8@380_d N_OUT7_Mp8@380_g N_VDD_Mp8@380_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@379 N_OUT8_Mn8@379_d N_OUT7_Mn8@379_g N_VSS_Mn8@379_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@378 N_OUT8_Mn8@378_d N_OUT7_Mn8@378_g N_VSS_Mn8@378_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@379 N_OUT8_Mp8@379_d N_OUT7_Mp8@379_g N_VDD_Mp8@379_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@378 N_OUT8_Mp8@378_d N_OUT7_Mp8@378_g N_VDD_Mp8@378_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@377 N_OUT8_Mn8@377_d N_OUT7_Mn8@377_g N_VSS_Mn8@377_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@376 N_OUT8_Mn8@376_d N_OUT7_Mn8@376_g N_VSS_Mn8@376_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@377 N_OUT8_Mp8@377_d N_OUT7_Mp8@377_g N_VDD_Mp8@377_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@376 N_OUT8_Mp8@376_d N_OUT7_Mp8@376_g N_VDD_Mp8@376_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@375 N_OUT8_Mn8@375_d N_OUT7_Mn8@375_g N_VSS_Mn8@375_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@374 N_OUT8_Mn8@374_d N_OUT7_Mn8@374_g N_VSS_Mn8@374_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@375 N_OUT8_Mp8@375_d N_OUT7_Mp8@375_g N_VDD_Mp8@375_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@374 N_OUT8_Mp8@374_d N_OUT7_Mp8@374_g N_VDD_Mp8@374_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@373 N_OUT8_Mn8@373_d N_OUT7_Mn8@373_g N_VSS_Mn8@373_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@372 N_OUT8_Mn8@372_d N_OUT7_Mn8@372_g N_VSS_Mn8@372_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@373 N_OUT8_Mp8@373_d N_OUT7_Mp8@373_g N_VDD_Mp8@373_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@372 N_OUT8_Mp8@372_d N_OUT7_Mp8@372_g N_VDD_Mp8@372_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@371 N_OUT8_Mn8@371_d N_OUT7_Mn8@371_g N_VSS_Mn8@371_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@370 N_OUT8_Mn8@370_d N_OUT7_Mn8@370_g N_VSS_Mn8@370_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@371 N_OUT8_Mp8@371_d N_OUT7_Mp8@371_g N_VDD_Mp8@371_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@370 N_OUT8_Mp8@370_d N_OUT7_Mp8@370_g N_VDD_Mp8@370_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@369 N_OUT8_Mn8@369_d N_OUT7_Mn8@369_g N_VSS_Mn8@369_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@368 N_OUT8_Mn8@368_d N_OUT7_Mn8@368_g N_VSS_Mn8@368_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@369 N_OUT8_Mp8@369_d N_OUT7_Mp8@369_g N_VDD_Mp8@369_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@368 N_OUT8_Mp8@368_d N_OUT7_Mp8@368_g N_VDD_Mp8@368_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@367 N_OUT8_Mn8@367_d N_OUT7_Mn8@367_g N_VSS_Mn8@367_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@366 N_OUT8_Mn8@366_d N_OUT7_Mn8@366_g N_VSS_Mn8@366_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@367 N_OUT8_Mp8@367_d N_OUT7_Mp8@367_g N_VDD_Mp8@367_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@366 N_OUT8_Mp8@366_d N_OUT7_Mp8@366_g N_VDD_Mp8@366_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@365 N_OUT8_Mn8@365_d N_OUT7_Mn8@365_g N_VSS_Mn8@365_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@364 N_OUT8_Mn8@364_d N_OUT7_Mn8@364_g N_VSS_Mn8@364_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@365 N_OUT8_Mp8@365_d N_OUT7_Mp8@365_g N_VDD_Mp8@365_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@364 N_OUT8_Mp8@364_d N_OUT7_Mp8@364_g N_VDD_Mp8@364_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@363 N_OUT8_Mn8@363_d N_OUT7_Mn8@363_g N_VSS_Mn8@363_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@362 N_OUT8_Mn8@362_d N_OUT7_Mn8@362_g N_VSS_Mn8@362_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@363 N_OUT8_Mp8@363_d N_OUT7_Mp8@363_g N_VDD_Mp8@363_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@362 N_OUT8_Mp8@362_d N_OUT7_Mp8@362_g N_VDD_Mp8@362_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@361 N_OUT8_Mn8@361_d N_OUT7_Mn8@361_g N_VSS_Mn8@361_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@360 N_OUT8_Mn8@360_d N_OUT7_Mn8@360_g N_VSS_Mn8@360_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@361 N_OUT8_Mp8@361_d N_OUT7_Mp8@361_g N_VDD_Mp8@361_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@360 N_OUT8_Mp8@360_d N_OUT7_Mp8@360_g N_VDD_Mp8@360_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@359 N_OUT8_Mn8@359_d N_OUT7_Mn8@359_g N_VSS_Mn8@359_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@358 N_OUT8_Mn8@358_d N_OUT7_Mn8@358_g N_VSS_Mn8@358_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@359 N_OUT8_Mp8@359_d N_OUT7_Mp8@359_g N_VDD_Mp8@359_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@358 N_OUT8_Mp8@358_d N_OUT7_Mp8@358_g N_VDD_Mp8@358_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@357 N_OUT8_Mn8@357_d N_OUT7_Mn8@357_g N_VSS_Mn8@357_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@356 N_OUT8_Mn8@356_d N_OUT7_Mn8@356_g N_VSS_Mn8@356_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@357 N_OUT8_Mp8@357_d N_OUT7_Mp8@357_g N_VDD_Mp8@357_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@356 N_OUT8_Mp8@356_d N_OUT7_Mp8@356_g N_VDD_Mp8@356_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@355 N_OUT8_Mn8@355_d N_OUT7_Mn8@355_g N_VSS_Mn8@355_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@354 N_OUT8_Mn8@354_d N_OUT7_Mn8@354_g N_VSS_Mn8@354_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@355 N_OUT8_Mp8@355_d N_OUT7_Mp8@355_g N_VDD_Mp8@355_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@354 N_OUT8_Mp8@354_d N_OUT7_Mp8@354_g N_VDD_Mp8@354_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@353 N_OUT8_Mn8@353_d N_OUT7_Mn8@353_g N_VSS_Mn8@353_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@352 N_OUT8_Mn8@352_d N_OUT7_Mn8@352_g N_VSS_Mn8@352_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@353 N_OUT8_Mp8@353_d N_OUT7_Mp8@353_g N_VDD_Mp8@353_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@352 N_OUT8_Mp8@352_d N_OUT7_Mp8@352_g N_VDD_Mp8@352_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@351 N_OUT8_Mn8@351_d N_OUT7_Mn8@351_g N_VSS_Mn8@351_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@350 N_OUT8_Mn8@350_d N_OUT7_Mn8@350_g N_VSS_Mn8@350_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@351 N_OUT8_Mp8@351_d N_OUT7_Mp8@351_g N_VDD_Mp8@351_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@350 N_OUT8_Mp8@350_d N_OUT7_Mp8@350_g N_VDD_Mp8@350_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@349 N_OUT8_Mn8@349_d N_OUT7_Mn8@349_g N_VSS_Mn8@349_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@348 N_OUT8_Mn8@348_d N_OUT7_Mn8@348_g N_VSS_Mn8@348_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@349 N_OUT8_Mp8@349_d N_OUT7_Mp8@349_g N_VDD_Mp8@349_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@348 N_OUT8_Mp8@348_d N_OUT7_Mp8@348_g N_VDD_Mp8@348_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@347 N_OUT8_Mn8@347_d N_OUT7_Mn8@347_g N_VSS_Mn8@347_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@346 N_OUT8_Mn8@346_d N_OUT7_Mn8@346_g N_VSS_Mn8@346_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@347 N_OUT8_Mp8@347_d N_OUT7_Mp8@347_g N_VDD_Mp8@347_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@346 N_OUT8_Mp8@346_d N_OUT7_Mp8@346_g N_VDD_Mp8@346_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@345 N_OUT8_Mn8@345_d N_OUT7_Mn8@345_g N_VSS_Mn8@345_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@344 N_OUT8_Mn8@344_d N_OUT7_Mn8@344_g N_VSS_Mn8@344_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@345 N_OUT8_Mp8@345_d N_OUT7_Mp8@345_g N_VDD_Mp8@345_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@344 N_OUT8_Mp8@344_d N_OUT7_Mp8@344_g N_VDD_Mp8@344_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@343 N_OUT8_Mn8@343_d N_OUT7_Mn8@343_g N_VSS_Mn8@343_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@342 N_OUT8_Mn8@342_d N_OUT7_Mn8@342_g N_VSS_Mn8@342_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@343 N_OUT8_Mp8@343_d N_OUT7_Mp8@343_g N_VDD_Mp8@343_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@342 N_OUT8_Mp8@342_d N_OUT7_Mp8@342_g N_VDD_Mp8@342_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@341 N_OUT8_Mn8@341_d N_OUT7_Mn8@341_g N_VSS_Mn8@341_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@340 N_OUT8_Mn8@340_d N_OUT7_Mn8@340_g N_VSS_Mn8@340_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@341 N_OUT8_Mp8@341_d N_OUT7_Mp8@341_g N_VDD_Mp8@341_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@340 N_OUT8_Mp8@340_d N_OUT7_Mp8@340_g N_VDD_Mp8@340_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@339 N_OUT8_Mn8@339_d N_OUT7_Mn8@339_g N_VSS_Mn8@339_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@338 N_OUT8_Mn8@338_d N_OUT7_Mn8@338_g N_VSS_Mn8@338_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@339 N_OUT8_Mp8@339_d N_OUT7_Mp8@339_g N_VDD_Mp8@339_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@338 N_OUT8_Mp8@338_d N_OUT7_Mp8@338_g N_VDD_Mp8@338_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@337 N_OUT8_Mn8@337_d N_OUT7_Mn8@337_g N_VSS_Mn8@337_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@336 N_OUT8_Mn8@336_d N_OUT7_Mn8@336_g N_VSS_Mn8@336_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@337 N_OUT8_Mp8@337_d N_OUT7_Mp8@337_g N_VDD_Mp8@337_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@336 N_OUT8_Mp8@336_d N_OUT7_Mp8@336_g N_VDD_Mp8@336_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@335 N_OUT8_Mn8@335_d N_OUT7_Mn8@335_g N_VSS_Mn8@335_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@334 N_OUT8_Mn8@334_d N_OUT7_Mn8@334_g N_VSS_Mn8@334_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@335 N_OUT8_Mp8@335_d N_OUT7_Mp8@335_g N_VDD_Mp8@335_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@334 N_OUT8_Mp8@334_d N_OUT7_Mp8@334_g N_VDD_Mp8@334_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@333 N_OUT8_Mn8@333_d N_OUT7_Mn8@333_g N_VSS_Mn8@333_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@332 N_OUT8_Mn8@332_d N_OUT7_Mn8@332_g N_VSS_Mn8@332_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@333 N_OUT8_Mp8@333_d N_OUT7_Mp8@333_g N_VDD_Mp8@333_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@332 N_OUT8_Mp8@332_d N_OUT7_Mp8@332_g N_VDD_Mp8@332_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@331 N_OUT8_Mn8@331_d N_OUT7_Mn8@331_g N_VSS_Mn8@331_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@330 N_OUT8_Mn8@330_d N_OUT7_Mn8@330_g N_VSS_Mn8@330_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@331 N_OUT8_Mp8@331_d N_OUT7_Mp8@331_g N_VDD_Mp8@331_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@330 N_OUT8_Mp8@330_d N_OUT7_Mp8@330_g N_VDD_Mp8@330_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@329 N_OUT8_Mn8@329_d N_OUT7_Mn8@329_g N_VSS_Mn8@329_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@328 N_OUT8_Mn8@328_d N_OUT7_Mn8@328_g N_VSS_Mn8@328_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@329 N_OUT8_Mp8@329_d N_OUT7_Mp8@329_g N_VDD_Mp8@329_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@328 N_OUT8_Mp8@328_d N_OUT7_Mp8@328_g N_VDD_Mp8@328_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@327 N_OUT8_Mn8@327_d N_OUT7_Mn8@327_g N_VSS_Mn8@327_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@326 N_OUT8_Mn8@326_d N_OUT7_Mn8@326_g N_VSS_Mn8@326_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@327 N_OUT8_Mp8@327_d N_OUT7_Mp8@327_g N_VDD_Mp8@327_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@326 N_OUT8_Mp8@326_d N_OUT7_Mp8@326_g N_VDD_Mp8@326_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@325 N_OUT8_Mn8@325_d N_OUT7_Mn8@325_g N_VSS_Mn8@325_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@324 N_OUT8_Mn8@324_d N_OUT7_Mn8@324_g N_VSS_Mn8@324_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@325 N_OUT8_Mp8@325_d N_OUT7_Mp8@325_g N_VDD_Mp8@325_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@324 N_OUT8_Mp8@324_d N_OUT7_Mp8@324_g N_VDD_Mp8@324_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@323 N_OUT8_Mn8@323_d N_OUT7_Mn8@323_g N_VSS_Mn8@323_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@322 N_OUT8_Mn8@322_d N_OUT7_Mn8@322_g N_VSS_Mn8@322_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@323 N_OUT8_Mp8@323_d N_OUT7_Mp8@323_g N_VDD_Mp8@323_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@322 N_OUT8_Mp8@322_d N_OUT7_Mp8@322_g N_VDD_Mp8@322_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@321 N_OUT8_Mn8@321_d N_OUT7_Mn8@321_g N_VSS_Mn8@321_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@320 N_OUT8_Mn8@320_d N_OUT7_Mn8@320_g N_VSS_Mn8@320_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@321 N_OUT8_Mp8@321_d N_OUT7_Mp8@321_g N_VDD_Mp8@321_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@320 N_OUT8_Mp8@320_d N_OUT7_Mp8@320_g N_VDD_Mp8@320_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@319 N_OUT8_Mn8@319_d N_OUT7_Mn8@319_g N_VSS_Mn8@319_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@318 N_OUT8_Mn8@318_d N_OUT7_Mn8@318_g N_VSS_Mn8@318_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@319 N_OUT8_Mp8@319_d N_OUT7_Mp8@319_g N_VDD_Mp8@319_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@318 N_OUT8_Mp8@318_d N_OUT7_Mp8@318_g N_VDD_Mp8@318_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@317 N_OUT8_Mn8@317_d N_OUT7_Mn8@317_g N_VSS_Mn8@317_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@316 N_OUT8_Mn8@316_d N_OUT7_Mn8@316_g N_VSS_Mn8@316_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@317 N_OUT8_Mp8@317_d N_OUT7_Mp8@317_g N_VDD_Mp8@317_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@316 N_OUT8_Mp8@316_d N_OUT7_Mp8@316_g N_VDD_Mp8@316_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@315 N_OUT8_Mn8@315_d N_OUT7_Mn8@315_g N_VSS_Mn8@315_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@314 N_OUT8_Mn8@314_d N_OUT7_Mn8@314_g N_VSS_Mn8@314_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@315 N_OUT8_Mp8@315_d N_OUT7_Mp8@315_g N_VDD_Mp8@315_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@314 N_OUT8_Mp8@314_d N_OUT7_Mp8@314_g N_VDD_Mp8@314_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@313 N_OUT8_Mn8@313_d N_OUT7_Mn8@313_g N_VSS_Mn8@313_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@312 N_OUT8_Mn8@312_d N_OUT7_Mn8@312_g N_VSS_Mn8@312_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@313 N_OUT8_Mp8@313_d N_OUT7_Mp8@313_g N_VDD_Mp8@313_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@312 N_OUT8_Mp8@312_d N_OUT7_Mp8@312_g N_VDD_Mp8@312_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@311 N_OUT8_Mn8@311_d N_OUT7_Mn8@311_g N_VSS_Mn8@311_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@310 N_OUT8_Mn8@310_d N_OUT7_Mn8@310_g N_VSS_Mn8@310_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@311 N_OUT8_Mp8@311_d N_OUT7_Mp8@311_g N_VDD_Mp8@311_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@310 N_OUT8_Mp8@310_d N_OUT7_Mp8@310_g N_VDD_Mp8@310_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@309 N_OUT8_Mn8@309_d N_OUT7_Mn8@309_g N_VSS_Mn8@309_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@308 N_OUT8_Mn8@308_d N_OUT7_Mn8@308_g N_VSS_Mn8@308_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@309 N_OUT8_Mp8@309_d N_OUT7_Mp8@309_g N_VDD_Mp8@309_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@308 N_OUT8_Mp8@308_d N_OUT7_Mp8@308_g N_VDD_Mp8@308_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@307 N_OUT8_Mn8@307_d N_OUT7_Mn8@307_g N_VSS_Mn8@307_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@306 N_OUT8_Mn8@306_d N_OUT7_Mn8@306_g N_VSS_Mn8@306_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@307 N_OUT8_Mp8@307_d N_OUT7_Mp8@307_g N_VDD_Mp8@307_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@306 N_OUT8_Mp8@306_d N_OUT7_Mp8@306_g N_VDD_Mp8@306_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@305 N_OUT8_Mn8@305_d N_OUT7_Mn8@305_g N_VSS_Mn8@305_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@304 N_OUT8_Mn8@304_d N_OUT7_Mn8@304_g N_VSS_Mn8@304_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@305 N_OUT8_Mp8@305_d N_OUT7_Mp8@305_g N_VDD_Mp8@305_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@304 N_OUT8_Mp8@304_d N_OUT7_Mp8@304_g N_VDD_Mp8@304_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@303 N_OUT8_Mn8@303_d N_OUT7_Mn8@303_g N_VSS_Mn8@303_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@302 N_OUT8_Mn8@302_d N_OUT7_Mn8@302_g N_VSS_Mn8@302_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@303 N_OUT8_Mp8@303_d N_OUT7_Mp8@303_g N_VDD_Mp8@303_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@302 N_OUT8_Mp8@302_d N_OUT7_Mp8@302_g N_VDD_Mp8@302_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@301 N_OUT8_Mn8@301_d N_OUT7_Mn8@301_g N_VSS_Mn8@301_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@300 N_OUT8_Mn8@300_d N_OUT7_Mn8@300_g N_VSS_Mn8@300_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@301 N_OUT8_Mp8@301_d N_OUT7_Mp8@301_g N_VDD_Mp8@301_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@300 N_OUT8_Mp8@300_d N_OUT7_Mp8@300_g N_VDD_Mp8@300_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@299 N_OUT8_Mn8@299_d N_OUT7_Mn8@299_g N_VSS_Mn8@299_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@298 N_OUT8_Mn8@298_d N_OUT7_Mn8@298_g N_VSS_Mn8@298_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@299 N_OUT8_Mp8@299_d N_OUT7_Mp8@299_g N_VDD_Mp8@299_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@298 N_OUT8_Mp8@298_d N_OUT7_Mp8@298_g N_VDD_Mp8@298_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@297 N_OUT8_Mn8@297_d N_OUT7_Mn8@297_g N_VSS_Mn8@297_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@296 N_OUT8_Mn8@296_d N_OUT7_Mn8@296_g N_VSS_Mn8@296_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@297 N_OUT8_Mp8@297_d N_OUT7_Mp8@297_g N_VDD_Mp8@297_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@296 N_OUT8_Mp8@296_d N_OUT7_Mp8@296_g N_VDD_Mp8@296_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@295 N_OUT8_Mn8@295_d N_OUT7_Mn8@295_g N_VSS_Mn8@295_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@294 N_OUT8_Mn8@294_d N_OUT7_Mn8@294_g N_VSS_Mn8@294_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@295 N_OUT8_Mp8@295_d N_OUT7_Mp8@295_g N_VDD_Mp8@295_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@294 N_OUT8_Mp8@294_d N_OUT7_Mp8@294_g N_VDD_Mp8@294_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@293 N_OUT8_Mn8@293_d N_OUT7_Mn8@293_g N_VSS_Mn8@293_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@292 N_OUT8_Mn8@292_d N_OUT7_Mn8@292_g N_VSS_Mn8@292_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@293 N_OUT8_Mp8@293_d N_OUT7_Mp8@293_g N_VDD_Mp8@293_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@292 N_OUT8_Mp8@292_d N_OUT7_Mp8@292_g N_VDD_Mp8@292_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@291 N_OUT8_Mn8@291_d N_OUT7_Mn8@291_g N_VSS_Mn8@291_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@290 N_OUT8_Mn8@290_d N_OUT7_Mn8@290_g N_VSS_Mn8@290_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@291 N_OUT8_Mp8@291_d N_OUT7_Mp8@291_g N_VDD_Mp8@291_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@290 N_OUT8_Mp8@290_d N_OUT7_Mp8@290_g N_VDD_Mp8@290_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@289 N_OUT8_Mn8@289_d N_OUT7_Mn8@289_g N_VSS_Mn8@289_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@288 N_OUT8_Mn8@288_d N_OUT7_Mn8@288_g N_VSS_Mn8@288_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@289 N_OUT8_Mp8@289_d N_OUT7_Mp8@289_g N_VDD_Mp8@289_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@288 N_OUT8_Mp8@288_d N_OUT7_Mp8@288_g N_VDD_Mp8@288_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@287 N_OUT8_Mn8@287_d N_OUT7_Mn8@287_g N_VSS_Mn8@287_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@286 N_OUT8_Mn8@286_d N_OUT7_Mn8@286_g N_VSS_Mn8@286_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@287 N_OUT8_Mp8@287_d N_OUT7_Mp8@287_g N_VDD_Mp8@287_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@286 N_OUT8_Mp8@286_d N_OUT7_Mp8@286_g N_VDD_Mp8@286_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@285 N_OUT8_Mn8@285_d N_OUT7_Mn8@285_g N_VSS_Mn8@285_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@284 N_OUT8_Mn8@284_d N_OUT7_Mn8@284_g N_VSS_Mn8@284_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@285 N_OUT8_Mp8@285_d N_OUT7_Mp8@285_g N_VDD_Mp8@285_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@284 N_OUT8_Mp8@284_d N_OUT7_Mp8@284_g N_VDD_Mp8@284_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@283 N_OUT8_Mn8@283_d N_OUT7_Mn8@283_g N_VSS_Mn8@283_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@282 N_OUT8_Mn8@282_d N_OUT7_Mn8@282_g N_VSS_Mn8@282_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@283 N_OUT8_Mp8@283_d N_OUT7_Mp8@283_g N_VDD_Mp8@283_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@282 N_OUT8_Mp8@282_d N_OUT7_Mp8@282_g N_VDD_Mp8@282_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@281 N_OUT8_Mn8@281_d N_OUT7_Mn8@281_g N_VSS_Mn8@281_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@280 N_OUT8_Mn8@280_d N_OUT7_Mn8@280_g N_VSS_Mn8@280_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@281 N_OUT8_Mp8@281_d N_OUT7_Mp8@281_g N_VDD_Mp8@281_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@280 N_OUT8_Mp8@280_d N_OUT7_Mp8@280_g N_VDD_Mp8@280_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@279 N_OUT8_Mn8@279_d N_OUT7_Mn8@279_g N_VSS_Mn8@279_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@278 N_OUT8_Mn8@278_d N_OUT7_Mn8@278_g N_VSS_Mn8@278_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@279 N_OUT8_Mp8@279_d N_OUT7_Mp8@279_g N_VDD_Mp8@279_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@278 N_OUT8_Mp8@278_d N_OUT7_Mp8@278_g N_VDD_Mp8@278_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@277 N_OUT8_Mn8@277_d N_OUT7_Mn8@277_g N_VSS_Mn8@277_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@276 N_OUT8_Mn8@276_d N_OUT7_Mn8@276_g N_VSS_Mn8@276_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@277 N_OUT8_Mp8@277_d N_OUT7_Mp8@277_g N_VDD_Mp8@277_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@276 N_OUT8_Mp8@276_d N_OUT7_Mp8@276_g N_VDD_Mp8@276_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@275 N_OUT8_Mn8@275_d N_OUT7_Mn8@275_g N_VSS_Mn8@275_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@274 N_OUT8_Mn8@274_d N_OUT7_Mn8@274_g N_VSS_Mn8@274_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@275 N_OUT8_Mp8@275_d N_OUT7_Mp8@275_g N_VDD_Mp8@275_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@274 N_OUT8_Mp8@274_d N_OUT7_Mp8@274_g N_VDD_Mp8@274_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@273 N_OUT8_Mn8@273_d N_OUT7_Mn8@273_g N_VSS_Mn8@273_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@272 N_OUT8_Mn8@272_d N_OUT7_Mn8@272_g N_VSS_Mn8@272_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@273 N_OUT8_Mp8@273_d N_OUT7_Mp8@273_g N_VDD_Mp8@273_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@272 N_OUT8_Mp8@272_d N_OUT7_Mp8@272_g N_VDD_Mp8@272_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@271 N_OUT8_Mn8@271_d N_OUT7_Mn8@271_g N_VSS_Mn8@271_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@270 N_OUT8_Mn8@270_d N_OUT7_Mn8@270_g N_VSS_Mn8@270_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@271 N_OUT8_Mp8@271_d N_OUT7_Mp8@271_g N_VDD_Mp8@271_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@270 N_OUT8_Mp8@270_d N_OUT7_Mp8@270_g N_VDD_Mp8@270_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@269 N_OUT8_Mn8@269_d N_OUT7_Mn8@269_g N_VSS_Mn8@269_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@268 N_OUT8_Mn8@268_d N_OUT7_Mn8@268_g N_VSS_Mn8@268_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@269 N_OUT8_Mp8@269_d N_OUT7_Mp8@269_g N_VDD_Mp8@269_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@268 N_OUT8_Mp8@268_d N_OUT7_Mp8@268_g N_VDD_Mp8@268_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@267 N_OUT8_Mn8@267_d N_OUT7_Mn8@267_g N_VSS_Mn8@267_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@266 N_OUT8_Mn8@266_d N_OUT7_Mn8@266_g N_VSS_Mn8@266_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@267 N_OUT8_Mp8@267_d N_OUT7_Mp8@267_g N_VDD_Mp8@267_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@266 N_OUT8_Mp8@266_d N_OUT7_Mp8@266_g N_VDD_Mp8@266_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@265 N_OUT8_Mn8@265_d N_OUT7_Mn8@265_g N_VSS_Mn8@265_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@264 N_OUT8_Mn8@264_d N_OUT7_Mn8@264_g N_VSS_Mn8@264_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@265 N_OUT8_Mp8@265_d N_OUT7_Mp8@265_g N_VDD_Mp8@265_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@264 N_OUT8_Mp8@264_d N_OUT7_Mp8@264_g N_VDD_Mp8@264_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@263 N_OUT8_Mn8@263_d N_OUT7_Mn8@263_g N_VSS_Mn8@263_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@262 N_OUT8_Mn8@262_d N_OUT7_Mn8@262_g N_VSS_Mn8@262_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@263 N_OUT8_Mp8@263_d N_OUT7_Mp8@263_g N_VDD_Mp8@263_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@262 N_OUT8_Mp8@262_d N_OUT7_Mp8@262_g N_VDD_Mp8@262_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@261 N_OUT8_Mn8@261_d N_OUT7_Mn8@261_g N_VSS_Mn8@261_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@260 N_OUT8_Mn8@260_d N_OUT7_Mn8@260_g N_VSS_Mn8@260_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@261 N_OUT8_Mp8@261_d N_OUT7_Mp8@261_g N_VDD_Mp8@261_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@260 N_OUT8_Mp8@260_d N_OUT7_Mp8@260_g N_VDD_Mp8@260_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@259 N_OUT8_Mn8@259_d N_OUT7_Mn8@259_g N_VSS_Mn8@259_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@258 N_OUT8_Mn8@258_d N_OUT7_Mn8@258_g N_VSS_Mn8@258_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@259 N_OUT8_Mp8@259_d N_OUT7_Mp8@259_g N_VDD_Mp8@259_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@258 N_OUT8_Mp8@258_d N_OUT7_Mp8@258_g N_VDD_Mp8@258_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@257 N_OUT8_Mn8@257_d N_OUT7_Mn8@257_g N_VSS_Mn8@257_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@256 N_OUT8_Mn8@256_d N_OUT7_Mn8@256_g N_VSS_Mn8@256_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@257 N_OUT8_Mp8@257_d N_OUT7_Mp8@257_g N_VDD_Mp8@257_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@256 N_OUT8_Mp8@256_d N_OUT7_Mp8@256_g N_VDD_Mp8@256_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@255 N_OUT8_Mn8@255_d N_OUT7_Mn8@255_g N_VSS_Mn8@255_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@254 N_OUT8_Mn8@254_d N_OUT7_Mn8@254_g N_VSS_Mn8@254_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@255 N_OUT8_Mp8@255_d N_OUT7_Mp8@255_g N_VDD_Mp8@255_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@254 N_OUT8_Mp8@254_d N_OUT7_Mp8@254_g N_VDD_Mp8@254_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@253 N_OUT8_Mn8@253_d N_OUT7_Mn8@253_g N_VSS_Mn8@253_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@252 N_OUT8_Mn8@252_d N_OUT7_Mn8@252_g N_VSS_Mn8@252_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@253 N_OUT8_Mp8@253_d N_OUT7_Mp8@253_g N_VDD_Mp8@253_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@252 N_OUT8_Mp8@252_d N_OUT7_Mp8@252_g N_VDD_Mp8@252_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@251 N_OUT8_Mn8@251_d N_OUT7_Mn8@251_g N_VSS_Mn8@251_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@250 N_OUT8_Mn8@250_d N_OUT7_Mn8@250_g N_VSS_Mn8@250_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@251 N_OUT8_Mp8@251_d N_OUT7_Mp8@251_g N_VDD_Mp8@251_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@250 N_OUT8_Mp8@250_d N_OUT7_Mp8@250_g N_VDD_Mp8@250_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@249 N_OUT8_Mn8@249_d N_OUT7_Mn8@249_g N_VSS_Mn8@249_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@248 N_OUT8_Mn8@248_d N_OUT7_Mn8@248_g N_VSS_Mn8@248_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@249 N_OUT8_Mp8@249_d N_OUT7_Mp8@249_g N_VDD_Mp8@249_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@248 N_OUT8_Mp8@248_d N_OUT7_Mp8@248_g N_VDD_Mp8@248_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@247 N_OUT8_Mn8@247_d N_OUT7_Mn8@247_g N_VSS_Mn8@247_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@246 N_OUT8_Mn8@246_d N_OUT7_Mn8@246_g N_VSS_Mn8@246_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@247 N_OUT8_Mp8@247_d N_OUT7_Mp8@247_g N_VDD_Mp8@247_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@246 N_OUT8_Mp8@246_d N_OUT7_Mp8@246_g N_VDD_Mp8@246_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@245 N_OUT8_Mn8@245_d N_OUT7_Mn8@245_g N_VSS_Mn8@245_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@244 N_OUT8_Mn8@244_d N_OUT7_Mn8@244_g N_VSS_Mn8@244_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@245 N_OUT8_Mp8@245_d N_OUT7_Mp8@245_g N_VDD_Mp8@245_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@244 N_OUT8_Mp8@244_d N_OUT7_Mp8@244_g N_VDD_Mp8@244_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@243 N_OUT8_Mn8@243_d N_OUT7_Mn8@243_g N_VSS_Mn8@243_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@242 N_OUT8_Mn8@242_d N_OUT7_Mn8@242_g N_VSS_Mn8@242_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@243 N_OUT8_Mp8@243_d N_OUT7_Mp8@243_g N_VDD_Mp8@243_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@242 N_OUT8_Mp8@242_d N_OUT7_Mp8@242_g N_VDD_Mp8@242_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@241 N_OUT8_Mn8@241_d N_OUT7_Mn8@241_g N_VSS_Mn8@241_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@240 N_OUT8_Mn8@240_d N_OUT7_Mn8@240_g N_VSS_Mn8@240_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@241 N_OUT8_Mp8@241_d N_OUT7_Mp8@241_g N_VDD_Mp8@241_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@240 N_OUT8_Mp8@240_d N_OUT7_Mp8@240_g N_VDD_Mp8@240_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@239 N_OUT8_Mn8@239_d N_OUT7_Mn8@239_g N_VSS_Mn8@239_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@238 N_OUT8_Mn8@238_d N_OUT7_Mn8@238_g N_VSS_Mn8@238_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@239 N_OUT8_Mp8@239_d N_OUT7_Mp8@239_g N_VDD_Mp8@239_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@238 N_OUT8_Mp8@238_d N_OUT7_Mp8@238_g N_VDD_Mp8@238_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@237 N_OUT8_Mn8@237_d N_OUT7_Mn8@237_g N_VSS_Mn8@237_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@236 N_OUT8_Mn8@236_d N_OUT7_Mn8@236_g N_VSS_Mn8@236_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@237 N_OUT8_Mp8@237_d N_OUT7_Mp8@237_g N_VDD_Mp8@237_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@236 N_OUT8_Mp8@236_d N_OUT7_Mp8@236_g N_VDD_Mp8@236_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@235 N_OUT8_Mn8@235_d N_OUT7_Mn8@235_g N_VSS_Mn8@235_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@234 N_OUT8_Mn8@234_d N_OUT7_Mn8@234_g N_VSS_Mn8@234_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@235 N_OUT8_Mp8@235_d N_OUT7_Mp8@235_g N_VDD_Mp8@235_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@234 N_OUT8_Mp8@234_d N_OUT7_Mp8@234_g N_VDD_Mp8@234_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@233 N_OUT8_Mn8@233_d N_OUT7_Mn8@233_g N_VSS_Mn8@233_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@232 N_OUT8_Mn8@232_d N_OUT7_Mn8@232_g N_VSS_Mn8@232_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@233 N_OUT8_Mp8@233_d N_OUT7_Mp8@233_g N_VDD_Mp8@233_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@232 N_OUT8_Mp8@232_d N_OUT7_Mp8@232_g N_VDD_Mp8@232_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@231 N_OUT8_Mn8@231_d N_OUT7_Mn8@231_g N_VSS_Mn8@231_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@230 N_OUT8_Mn8@230_d N_OUT7_Mn8@230_g N_VSS_Mn8@230_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@231 N_OUT8_Mp8@231_d N_OUT7_Mp8@231_g N_VDD_Mp8@231_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@230 N_OUT8_Mp8@230_d N_OUT7_Mp8@230_g N_VDD_Mp8@230_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@229 N_OUT8_Mn8@229_d N_OUT7_Mn8@229_g N_VSS_Mn8@229_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@228 N_OUT8_Mn8@228_d N_OUT7_Mn8@228_g N_VSS_Mn8@228_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@229 N_OUT8_Mp8@229_d N_OUT7_Mp8@229_g N_VDD_Mp8@229_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@228 N_OUT8_Mp8@228_d N_OUT7_Mp8@228_g N_VDD_Mp8@228_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@227 N_OUT8_Mn8@227_d N_OUT7_Mn8@227_g N_VSS_Mn8@227_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@226 N_OUT8_Mn8@226_d N_OUT7_Mn8@226_g N_VSS_Mn8@226_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@227 N_OUT8_Mp8@227_d N_OUT7_Mp8@227_g N_VDD_Mp8@227_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@226 N_OUT8_Mp8@226_d N_OUT7_Mp8@226_g N_VDD_Mp8@226_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@225 N_OUT8_Mn8@225_d N_OUT7_Mn8@225_g N_VSS_Mn8@225_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@224 N_OUT8_Mn8@224_d N_OUT7_Mn8@224_g N_VSS_Mn8@224_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@225 N_OUT8_Mp8@225_d N_OUT7_Mp8@225_g N_VDD_Mp8@225_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@224 N_OUT8_Mp8@224_d N_OUT7_Mp8@224_g N_VDD_Mp8@224_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@223 N_OUT8_Mn8@223_d N_OUT7_Mn8@223_g N_VSS_Mn8@223_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@222 N_OUT8_Mn8@222_d N_OUT7_Mn8@222_g N_VSS_Mn8@222_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@223 N_OUT8_Mp8@223_d N_OUT7_Mp8@223_g N_VDD_Mp8@223_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@222 N_OUT8_Mp8@222_d N_OUT7_Mp8@222_g N_VDD_Mp8@222_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@221 N_OUT8_Mn8@221_d N_OUT7_Mn8@221_g N_VSS_Mn8@221_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@220 N_OUT8_Mn8@220_d N_OUT7_Mn8@220_g N_VSS_Mn8@220_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@221 N_OUT8_Mp8@221_d N_OUT7_Mp8@221_g N_VDD_Mp8@221_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@220 N_OUT8_Mp8@220_d N_OUT7_Mp8@220_g N_VDD_Mp8@220_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@219 N_OUT8_Mn8@219_d N_OUT7_Mn8@219_g N_VSS_Mn8@219_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@218 N_OUT8_Mn8@218_d N_OUT7_Mn8@218_g N_VSS_Mn8@218_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@219 N_OUT8_Mp8@219_d N_OUT7_Mp8@219_g N_VDD_Mp8@219_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@218 N_OUT8_Mp8@218_d N_OUT7_Mp8@218_g N_VDD_Mp8@218_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@217 N_OUT8_Mn8@217_d N_OUT7_Mn8@217_g N_VSS_Mn8@217_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@216 N_OUT8_Mn8@216_d N_OUT7_Mn8@216_g N_VSS_Mn8@216_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@217 N_OUT8_Mp8@217_d N_OUT7_Mp8@217_g N_VDD_Mp8@217_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@216 N_OUT8_Mp8@216_d N_OUT7_Mp8@216_g N_VDD_Mp8@216_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@215 N_OUT8_Mn8@215_d N_OUT7_Mn8@215_g N_VSS_Mn8@215_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@214 N_OUT8_Mn8@214_d N_OUT7_Mn8@214_g N_VSS_Mn8@214_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@215 N_OUT8_Mp8@215_d N_OUT7_Mp8@215_g N_VDD_Mp8@215_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@214 N_OUT8_Mp8@214_d N_OUT7_Mp8@214_g N_VDD_Mp8@214_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@213 N_OUT8_Mn8@213_d N_OUT7_Mn8@213_g N_VSS_Mn8@213_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@212 N_OUT8_Mn8@212_d N_OUT7_Mn8@212_g N_VSS_Mn8@212_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@213 N_OUT8_Mp8@213_d N_OUT7_Mp8@213_g N_VDD_Mp8@213_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@212 N_OUT8_Mp8@212_d N_OUT7_Mp8@212_g N_VDD_Mp8@212_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@211 N_OUT8_Mn8@211_d N_OUT7_Mn8@211_g N_VSS_Mn8@211_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@210 N_OUT8_Mn8@210_d N_OUT7_Mn8@210_g N_VSS_Mn8@210_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@211 N_OUT8_Mp8@211_d N_OUT7_Mp8@211_g N_VDD_Mp8@211_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@210 N_OUT8_Mp8@210_d N_OUT7_Mp8@210_g N_VDD_Mp8@210_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@209 N_OUT8_Mn8@209_d N_OUT7_Mn8@209_g N_VSS_Mn8@209_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@208 N_OUT8_Mn8@208_d N_OUT7_Mn8@208_g N_VSS_Mn8@208_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@209 N_OUT8_Mp8@209_d N_OUT7_Mp8@209_g N_VDD_Mp8@209_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@208 N_OUT8_Mp8@208_d N_OUT7_Mp8@208_g N_VDD_Mp8@208_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@207 N_OUT8_Mn8@207_d N_OUT7_Mn8@207_g N_VSS_Mn8@207_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@206 N_OUT8_Mn8@206_d N_OUT7_Mn8@206_g N_VSS_Mn8@206_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@207 N_OUT8_Mp8@207_d N_OUT7_Mp8@207_g N_VDD_Mp8@207_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@206 N_OUT8_Mp8@206_d N_OUT7_Mp8@206_g N_VDD_Mp8@206_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@205 N_OUT8_Mn8@205_d N_OUT7_Mn8@205_g N_VSS_Mn8@205_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@204 N_OUT8_Mn8@204_d N_OUT7_Mn8@204_g N_VSS_Mn8@204_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@205 N_OUT8_Mp8@205_d N_OUT7_Mp8@205_g N_VDD_Mp8@205_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@204 N_OUT8_Mp8@204_d N_OUT7_Mp8@204_g N_VDD_Mp8@204_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@203 N_OUT8_Mn8@203_d N_OUT7_Mn8@203_g N_VSS_Mn8@203_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@202 N_OUT8_Mn8@202_d N_OUT7_Mn8@202_g N_VSS_Mn8@202_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@203 N_OUT8_Mp8@203_d N_OUT7_Mp8@203_g N_VDD_Mp8@203_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@202 N_OUT8_Mp8@202_d N_OUT7_Mp8@202_g N_VDD_Mp8@202_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@201 N_OUT8_Mn8@201_d N_OUT7_Mn8@201_g N_VSS_Mn8@201_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@200 N_OUT8_Mn8@200_d N_OUT7_Mn8@200_g N_VSS_Mn8@200_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@201 N_OUT8_Mp8@201_d N_OUT7_Mp8@201_g N_VDD_Mp8@201_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@200 N_OUT8_Mp8@200_d N_OUT7_Mp8@200_g N_VDD_Mp8@200_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@199 N_OUT8_Mn8@199_d N_OUT7_Mn8@199_g N_VSS_Mn8@199_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@198 N_OUT8_Mn8@198_d N_OUT7_Mn8@198_g N_VSS_Mn8@198_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@199 N_OUT8_Mp8@199_d N_OUT7_Mp8@199_g N_VDD_Mp8@199_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@198 N_OUT8_Mp8@198_d N_OUT7_Mp8@198_g N_VDD_Mp8@198_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@197 N_OUT8_Mn8@197_d N_OUT7_Mn8@197_g N_VSS_Mn8@197_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@196 N_OUT8_Mn8@196_d N_OUT7_Mn8@196_g N_VSS_Mn8@196_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@197 N_OUT8_Mp8@197_d N_OUT7_Mp8@197_g N_VDD_Mp8@197_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@196 N_OUT8_Mp8@196_d N_OUT7_Mp8@196_g N_VDD_Mp8@196_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@195 N_OUT8_Mn8@195_d N_OUT7_Mn8@195_g N_VSS_Mn8@195_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@194 N_OUT8_Mn8@194_d N_OUT7_Mn8@194_g N_VSS_Mn8@194_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@195 N_OUT8_Mp8@195_d N_OUT7_Mp8@195_g N_VDD_Mp8@195_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@194 N_OUT8_Mp8@194_d N_OUT7_Mp8@194_g N_VDD_Mp8@194_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@193 N_OUT8_Mn8@193_d N_OUT7_Mn8@193_g N_VSS_Mn8@193_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@192 N_OUT8_Mn8@192_d N_OUT7_Mn8@192_g N_VSS_Mn8@192_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@193 N_OUT8_Mp8@193_d N_OUT7_Mp8@193_g N_VDD_Mp8@193_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@192 N_OUT8_Mp8@192_d N_OUT7_Mp8@192_g N_VDD_Mp8@192_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@191 N_OUT8_Mn8@191_d N_OUT7_Mn8@191_g N_VSS_Mn8@191_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@190 N_OUT8_Mn8@190_d N_OUT7_Mn8@190_g N_VSS_Mn8@190_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@191 N_OUT8_Mp8@191_d N_OUT7_Mp8@191_g N_VDD_Mp8@191_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@190 N_OUT8_Mp8@190_d N_OUT7_Mp8@190_g N_VDD_Mp8@190_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@189 N_OUT8_Mn8@189_d N_OUT7_Mn8@189_g N_VSS_Mn8@189_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@188 N_OUT8_Mn8@188_d N_OUT7_Mn8@188_g N_VSS_Mn8@188_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@189 N_OUT8_Mp8@189_d N_OUT7_Mp8@189_g N_VDD_Mp8@189_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@188 N_OUT8_Mp8@188_d N_OUT7_Mp8@188_g N_VDD_Mp8@188_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@187 N_OUT8_Mn8@187_d N_OUT7_Mn8@187_g N_VSS_Mn8@187_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@186 N_OUT8_Mn8@186_d N_OUT7_Mn8@186_g N_VSS_Mn8@186_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@187 N_OUT8_Mp8@187_d N_OUT7_Mp8@187_g N_VDD_Mp8@187_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@186 N_OUT8_Mp8@186_d N_OUT7_Mp8@186_g N_VDD_Mp8@186_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@185 N_OUT8_Mn8@185_d N_OUT7_Mn8@185_g N_VSS_Mn8@185_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@184 N_OUT8_Mn8@184_d N_OUT7_Mn8@184_g N_VSS_Mn8@184_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@185 N_OUT8_Mp8@185_d N_OUT7_Mp8@185_g N_VDD_Mp8@185_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@184 N_OUT8_Mp8@184_d N_OUT7_Mp8@184_g N_VDD_Mp8@184_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@183 N_OUT8_Mn8@183_d N_OUT7_Mn8@183_g N_VSS_Mn8@183_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@182 N_OUT8_Mn8@182_d N_OUT7_Mn8@182_g N_VSS_Mn8@182_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@183 N_OUT8_Mp8@183_d N_OUT7_Mp8@183_g N_VDD_Mp8@183_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@182 N_OUT8_Mp8@182_d N_OUT7_Mp8@182_g N_VDD_Mp8@182_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@181 N_OUT8_Mn8@181_d N_OUT7_Mn8@181_g N_VSS_Mn8@181_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@180 N_OUT8_Mn8@180_d N_OUT7_Mn8@180_g N_VSS_Mn8@180_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@181 N_OUT8_Mp8@181_d N_OUT7_Mp8@181_g N_VDD_Mp8@181_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@180 N_OUT8_Mp8@180_d N_OUT7_Mp8@180_g N_VDD_Mp8@180_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@179 N_OUT8_Mn8@179_d N_OUT7_Mn8@179_g N_VSS_Mn8@179_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@178 N_OUT8_Mn8@178_d N_OUT7_Mn8@178_g N_VSS_Mn8@178_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@179 N_OUT8_Mp8@179_d N_OUT7_Mp8@179_g N_VDD_Mp8@179_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@178 N_OUT8_Mp8@178_d N_OUT7_Mp8@178_g N_VDD_Mp8@178_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@177 N_OUT8_Mn8@177_d N_OUT7_Mn8@177_g N_VSS_Mn8@177_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@176 N_OUT8_Mn8@176_d N_OUT7_Mn8@176_g N_VSS_Mn8@176_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@177 N_OUT8_Mp8@177_d N_OUT7_Mp8@177_g N_VDD_Mp8@177_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@176 N_OUT8_Mp8@176_d N_OUT7_Mp8@176_g N_VDD_Mp8@176_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@175 N_OUT8_Mn8@175_d N_OUT7_Mn8@175_g N_VSS_Mn8@175_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@174 N_OUT8_Mn8@174_d N_OUT7_Mn8@174_g N_VSS_Mn8@174_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@175 N_OUT8_Mp8@175_d N_OUT7_Mp8@175_g N_VDD_Mp8@175_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@174 N_OUT8_Mp8@174_d N_OUT7_Mp8@174_g N_VDD_Mp8@174_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@173 N_OUT8_Mn8@173_d N_OUT7_Mn8@173_g N_VSS_Mn8@173_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@172 N_OUT8_Mn8@172_d N_OUT7_Mn8@172_g N_VSS_Mn8@172_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@173 N_OUT8_Mp8@173_d N_OUT7_Mp8@173_g N_VDD_Mp8@173_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@172 N_OUT8_Mp8@172_d N_OUT7_Mp8@172_g N_VDD_Mp8@172_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@171 N_OUT8_Mn8@171_d N_OUT7_Mn8@171_g N_VSS_Mn8@171_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@170 N_OUT8_Mn8@170_d N_OUT7_Mn8@170_g N_VSS_Mn8@170_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@171 N_OUT8_Mp8@171_d N_OUT7_Mp8@171_g N_VDD_Mp8@171_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@170 N_OUT8_Mp8@170_d N_OUT7_Mp8@170_g N_VDD_Mp8@170_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@169 N_OUT8_Mn8@169_d N_OUT7_Mn8@169_g N_VSS_Mn8@169_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@168 N_OUT8_Mn8@168_d N_OUT7_Mn8@168_g N_VSS_Mn8@168_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@169 N_OUT8_Mp8@169_d N_OUT7_Mp8@169_g N_VDD_Mp8@169_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@168 N_OUT8_Mp8@168_d N_OUT7_Mp8@168_g N_VDD_Mp8@168_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@167 N_OUT8_Mn8@167_d N_OUT7_Mn8@167_g N_VSS_Mn8@167_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@166 N_OUT8_Mn8@166_d N_OUT7_Mn8@166_g N_VSS_Mn8@166_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@167 N_OUT8_Mp8@167_d N_OUT7_Mp8@167_g N_VDD_Mp8@167_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@166 N_OUT8_Mp8@166_d N_OUT7_Mp8@166_g N_VDD_Mp8@166_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@165 N_OUT8_Mn8@165_d N_OUT7_Mn8@165_g N_VSS_Mn8@165_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@164 N_OUT8_Mn8@164_d N_OUT7_Mn8@164_g N_VSS_Mn8@164_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@165 N_OUT8_Mp8@165_d N_OUT7_Mp8@165_g N_VDD_Mp8@165_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@164 N_OUT8_Mp8@164_d N_OUT7_Mp8@164_g N_VDD_Mp8@164_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@163 N_OUT8_Mn8@163_d N_OUT7_Mn8@163_g N_VSS_Mn8@163_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@162 N_OUT8_Mn8@162_d N_OUT7_Mn8@162_g N_VSS_Mn8@162_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@163 N_OUT8_Mp8@163_d N_OUT7_Mp8@163_g N_VDD_Mp8@163_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@162 N_OUT8_Mp8@162_d N_OUT7_Mp8@162_g N_VDD_Mp8@162_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@161 N_OUT8_Mn8@161_d N_OUT7_Mn8@161_g N_VSS_Mn8@161_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@160 N_OUT8_Mn8@160_d N_OUT7_Mn8@160_g N_VSS_Mn8@160_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@161 N_OUT8_Mp8@161_d N_OUT7_Mp8@161_g N_VDD_Mp8@161_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@160 N_OUT8_Mp8@160_d N_OUT7_Mp8@160_g N_VDD_Mp8@160_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@159 N_OUT8_Mn8@159_d N_OUT7_Mn8@159_g N_VSS_Mn8@159_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@158 N_OUT8_Mn8@158_d N_OUT7_Mn8@158_g N_VSS_Mn8@158_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@159 N_OUT8_Mp8@159_d N_OUT7_Mp8@159_g N_VDD_Mp8@159_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@158 N_OUT8_Mp8@158_d N_OUT7_Mp8@158_g N_VDD_Mp8@158_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@157 N_OUT8_Mn8@157_d N_OUT7_Mn8@157_g N_VSS_Mn8@157_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@156 N_OUT8_Mn8@156_d N_OUT7_Mn8@156_g N_VSS_Mn8@156_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@157 N_OUT8_Mp8@157_d N_OUT7_Mp8@157_g N_VDD_Mp8@157_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@156 N_OUT8_Mp8@156_d N_OUT7_Mp8@156_g N_VDD_Mp8@156_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@155 N_OUT8_Mn8@155_d N_OUT7_Mn8@155_g N_VSS_Mn8@155_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@154 N_OUT8_Mn8@154_d N_OUT7_Mn8@154_g N_VSS_Mn8@154_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@155 N_OUT8_Mp8@155_d N_OUT7_Mp8@155_g N_VDD_Mp8@155_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@154 N_OUT8_Mp8@154_d N_OUT7_Mp8@154_g N_VDD_Mp8@154_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@153 N_OUT8_Mn8@153_d N_OUT7_Mn8@153_g N_VSS_Mn8@153_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@152 N_OUT8_Mn8@152_d N_OUT7_Mn8@152_g N_VSS_Mn8@152_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@153 N_OUT8_Mp8@153_d N_OUT7_Mp8@153_g N_VDD_Mp8@153_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@152 N_OUT8_Mp8@152_d N_OUT7_Mp8@152_g N_VDD_Mp8@152_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@151 N_OUT8_Mn8@151_d N_OUT7_Mn8@151_g N_VSS_Mn8@151_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@150 N_OUT8_Mn8@150_d N_OUT7_Mn8@150_g N_VSS_Mn8@150_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@151 N_OUT8_Mp8@151_d N_OUT7_Mp8@151_g N_VDD_Mp8@151_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@150 N_OUT8_Mp8@150_d N_OUT7_Mp8@150_g N_VDD_Mp8@150_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@149 N_OUT8_Mn8@149_d N_OUT7_Mn8@149_g N_VSS_Mn8@149_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@148 N_OUT8_Mn8@148_d N_OUT7_Mn8@148_g N_VSS_Mn8@148_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@149 N_OUT8_Mp8@149_d N_OUT7_Mp8@149_g N_VDD_Mp8@149_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@148 N_OUT8_Mp8@148_d N_OUT7_Mp8@148_g N_VDD_Mp8@148_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@147 N_OUT8_Mn8@147_d N_OUT7_Mn8@147_g N_VSS_Mn8@147_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@146 N_OUT8_Mn8@146_d N_OUT7_Mn8@146_g N_VSS_Mn8@146_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@147 N_OUT8_Mp8@147_d N_OUT7_Mp8@147_g N_VDD_Mp8@147_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@146 N_OUT8_Mp8@146_d N_OUT7_Mp8@146_g N_VDD_Mp8@146_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@145 N_OUT8_Mn8@145_d N_OUT7_Mn8@145_g N_VSS_Mn8@145_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@144 N_OUT8_Mn8@144_d N_OUT7_Mn8@144_g N_VSS_Mn8@144_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@145 N_OUT8_Mp8@145_d N_OUT7_Mp8@145_g N_VDD_Mp8@145_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@144 N_OUT8_Mp8@144_d N_OUT7_Mp8@144_g N_VDD_Mp8@144_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@143 N_OUT8_Mn8@143_d N_OUT7_Mn8@143_g N_VSS_Mn8@143_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@142 N_OUT8_Mn8@142_d N_OUT7_Mn8@142_g N_VSS_Mn8@142_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@143 N_OUT8_Mp8@143_d N_OUT7_Mp8@143_g N_VDD_Mp8@143_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@142 N_OUT8_Mp8@142_d N_OUT7_Mp8@142_g N_VDD_Mp8@142_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@141 N_OUT8_Mn8@141_d N_OUT7_Mn8@141_g N_VSS_Mn8@141_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@140 N_OUT8_Mn8@140_d N_OUT7_Mn8@140_g N_VSS_Mn8@140_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@141 N_OUT8_Mp8@141_d N_OUT7_Mp8@141_g N_VDD_Mp8@141_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@140 N_OUT8_Mp8@140_d N_OUT7_Mp8@140_g N_VDD_Mp8@140_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@139 N_OUT8_Mn8@139_d N_OUT7_Mn8@139_g N_VSS_Mn8@139_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@138 N_OUT8_Mn8@138_d N_OUT7_Mn8@138_g N_VSS_Mn8@138_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@139 N_OUT8_Mp8@139_d N_OUT7_Mp8@139_g N_VDD_Mp8@139_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@138 N_OUT8_Mp8@138_d N_OUT7_Mp8@138_g N_VDD_Mp8@138_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@137 N_OUT8_Mn8@137_d N_OUT7_Mn8@137_g N_VSS_Mn8@137_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@136 N_OUT8_Mn8@136_d N_OUT7_Mn8@136_g N_VSS_Mn8@136_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@137 N_OUT8_Mp8@137_d N_OUT7_Mp8@137_g N_VDD_Mp8@137_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@136 N_OUT8_Mp8@136_d N_OUT7_Mp8@136_g N_VDD_Mp8@136_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@135 N_OUT8_Mn8@135_d N_OUT7_Mn8@135_g N_VSS_Mn8@135_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@134 N_OUT8_Mn8@134_d N_OUT7_Mn8@134_g N_VSS_Mn8@134_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@135 N_OUT8_Mp8@135_d N_OUT7_Mp8@135_g N_VDD_Mp8@135_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@134 N_OUT8_Mp8@134_d N_OUT7_Mp8@134_g N_VDD_Mp8@134_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@133 N_OUT8_Mn8@133_d N_OUT7_Mn8@133_g N_VSS_Mn8@133_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@132 N_OUT8_Mn8@132_d N_OUT7_Mn8@132_g N_VSS_Mn8@132_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@133 N_OUT8_Mp8@133_d N_OUT7_Mp8@133_g N_VDD_Mp8@133_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@132 N_OUT8_Mp8@132_d N_OUT7_Mp8@132_g N_VDD_Mp8@132_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@131 N_OUT8_Mn8@131_d N_OUT7_Mn8@131_g N_VSS_Mn8@131_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@130 N_OUT8_Mn8@130_d N_OUT7_Mn8@130_g N_VSS_Mn8@130_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@131 N_OUT8_Mp8@131_d N_OUT7_Mp8@131_g N_VDD_Mp8@131_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@130 N_OUT8_Mp8@130_d N_OUT7_Mp8@130_g N_VDD_Mp8@130_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@129 N_OUT8_Mn8@129_d N_OUT7_Mn8@129_g N_VSS_Mn8@129_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@128 N_OUT8_Mn8@128_d N_OUT7_Mn8@128_g N_VSS_Mn8@128_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@129 N_OUT8_Mp8@129_d N_OUT7_Mp8@129_g N_VDD_Mp8@129_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@128 N_OUT8_Mp8@128_d N_OUT7_Mp8@128_g N_VDD_Mp8@128_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@127 N_OUT8_Mn8@127_d N_OUT7_Mn8@127_g N_VSS_Mn8@127_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@126 N_OUT8_Mn8@126_d N_OUT7_Mn8@126_g N_VSS_Mn8@126_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@127 N_OUT8_Mp8@127_d N_OUT7_Mp8@127_g N_VDD_Mp8@127_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@126 N_OUT8_Mp8@126_d N_OUT7_Mp8@126_g N_VDD_Mp8@126_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@125 N_OUT8_Mn8@125_d N_OUT7_Mn8@125_g N_VSS_Mn8@125_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@124 N_OUT8_Mn8@124_d N_OUT7_Mn8@124_g N_VSS_Mn8@124_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@125 N_OUT8_Mp8@125_d N_OUT7_Mp8@125_g N_VDD_Mp8@125_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@124 N_OUT8_Mp8@124_d N_OUT7_Mp8@124_g N_VDD_Mp8@124_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@123 N_OUT8_Mn8@123_d N_OUT7_Mn8@123_g N_VSS_Mn8@123_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@122 N_OUT8_Mn8@122_d N_OUT7_Mn8@122_g N_VSS_Mn8@122_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@123 N_OUT8_Mp8@123_d N_OUT7_Mp8@123_g N_VDD_Mp8@123_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@122 N_OUT8_Mp8@122_d N_OUT7_Mp8@122_g N_VDD_Mp8@122_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@121 N_OUT8_Mn8@121_d N_OUT7_Mn8@121_g N_VSS_Mn8@121_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@120 N_OUT8_Mn8@120_d N_OUT7_Mn8@120_g N_VSS_Mn8@120_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@121 N_OUT8_Mp8@121_d N_OUT7_Mp8@121_g N_VDD_Mp8@121_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@120 N_OUT8_Mp8@120_d N_OUT7_Mp8@120_g N_VDD_Mp8@120_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@119 N_OUT8_Mn8@119_d N_OUT7_Mn8@119_g N_VSS_Mn8@119_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@118 N_OUT8_Mn8@118_d N_OUT7_Mn8@118_g N_VSS_Mn8@118_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@119 N_OUT8_Mp8@119_d N_OUT7_Mp8@119_g N_VDD_Mp8@119_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@118 N_OUT8_Mp8@118_d N_OUT7_Mp8@118_g N_VDD_Mp8@118_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@117 N_OUT8_Mn8@117_d N_OUT7_Mn8@117_g N_VSS_Mn8@117_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@116 N_OUT8_Mn8@116_d N_OUT7_Mn8@116_g N_VSS_Mn8@116_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@117 N_OUT8_Mp8@117_d N_OUT7_Mp8@117_g N_VDD_Mp8@117_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@116 N_OUT8_Mp8@116_d N_OUT7_Mp8@116_g N_VDD_Mp8@116_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@115 N_OUT8_Mn8@115_d N_OUT7_Mn8@115_g N_VSS_Mn8@115_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@114 N_OUT8_Mn8@114_d N_OUT7_Mn8@114_g N_VSS_Mn8@114_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@115 N_OUT8_Mp8@115_d N_OUT7_Mp8@115_g N_VDD_Mp8@115_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@114 N_OUT8_Mp8@114_d N_OUT7_Mp8@114_g N_VDD_Mp8@114_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@113 N_OUT8_Mn8@113_d N_OUT7_Mn8@113_g N_VSS_Mn8@113_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@112 N_OUT8_Mn8@112_d N_OUT7_Mn8@112_g N_VSS_Mn8@112_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@113 N_OUT8_Mp8@113_d N_OUT7_Mp8@113_g N_VDD_Mp8@113_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@112 N_OUT8_Mp8@112_d N_OUT7_Mp8@112_g N_VDD_Mp8@112_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@111 N_OUT8_Mn8@111_d N_OUT7_Mn8@111_g N_VSS_Mn8@111_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@110 N_OUT8_Mn8@110_d N_OUT7_Mn8@110_g N_VSS_Mn8@110_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@111 N_OUT8_Mp8@111_d N_OUT7_Mp8@111_g N_VDD_Mp8@111_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@110 N_OUT8_Mp8@110_d N_OUT7_Mp8@110_g N_VDD_Mp8@110_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@109 N_OUT8_Mn8@109_d N_OUT7_Mn8@109_g N_VSS_Mn8@109_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@108 N_OUT8_Mn8@108_d N_OUT7_Mn8@108_g N_VSS_Mn8@108_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@109 N_OUT8_Mp8@109_d N_OUT7_Mp8@109_g N_VDD_Mp8@109_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@108 N_OUT8_Mp8@108_d N_OUT7_Mp8@108_g N_VDD_Mp8@108_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@107 N_OUT8_Mn8@107_d N_OUT7_Mn8@107_g N_VSS_Mn8@107_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@106 N_OUT8_Mn8@106_d N_OUT7_Mn8@106_g N_VSS_Mn8@106_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@107 N_OUT8_Mp8@107_d N_OUT7_Mp8@107_g N_VDD_Mp8@107_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@106 N_OUT8_Mp8@106_d N_OUT7_Mp8@106_g N_VDD_Mp8@106_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@105 N_OUT8_Mn8@105_d N_OUT7_Mn8@105_g N_VSS_Mn8@105_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@104 N_OUT8_Mn8@104_d N_OUT7_Mn8@104_g N_VSS_Mn8@104_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@105 N_OUT8_Mp8@105_d N_OUT7_Mp8@105_g N_VDD_Mp8@105_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@104 N_OUT8_Mp8@104_d N_OUT7_Mp8@104_g N_VDD_Mp8@104_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@103 N_OUT8_Mn8@103_d N_OUT7_Mn8@103_g N_VSS_Mn8@103_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@102 N_OUT8_Mn8@102_d N_OUT7_Mn8@102_g N_VSS_Mn8@102_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@103 N_OUT8_Mp8@103_d N_OUT7_Mp8@103_g N_VDD_Mp8@103_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@102 N_OUT8_Mp8@102_d N_OUT7_Mp8@102_g N_VDD_Mp8@102_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@101 N_OUT8_Mn8@101_d N_OUT7_Mn8@101_g N_VSS_Mn8@101_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@100 N_OUT8_Mn8@100_d N_OUT7_Mn8@100_g N_VSS_Mn8@100_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@101 N_OUT8_Mp8@101_d N_OUT7_Mp8@101_g N_VDD_Mp8@101_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@100 N_OUT8_Mp8@100_d N_OUT7_Mp8@100_g N_VDD_Mp8@100_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@99 N_OUT8_Mn8@99_d N_OUT7_Mn8@99_g N_VSS_Mn8@99_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@98 N_OUT8_Mn8@98_d N_OUT7_Mn8@98_g N_VSS_Mn8@98_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@99 N_OUT8_Mp8@99_d N_OUT7_Mp8@99_g N_VDD_Mp8@99_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@98 N_OUT8_Mp8@98_d N_OUT7_Mp8@98_g N_VDD_Mp8@98_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@97 N_OUT8_Mn8@97_d N_OUT7_Mn8@97_g N_VSS_Mn8@97_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@96 N_OUT8_Mn8@96_d N_OUT7_Mn8@96_g N_VSS_Mn8@96_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@97 N_OUT8_Mp8@97_d N_OUT7_Mp8@97_g N_VDD_Mp8@97_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@96 N_OUT8_Mp8@96_d N_OUT7_Mp8@96_g N_VDD_Mp8@96_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@95 N_OUT8_Mn8@95_d N_OUT7_Mn8@95_g N_VSS_Mn8@95_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@94 N_OUT8_Mn8@94_d N_OUT7_Mn8@94_g N_VSS_Mn8@94_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@95 N_OUT8_Mp8@95_d N_OUT7_Mp8@95_g N_VDD_Mp8@95_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@94 N_OUT8_Mp8@94_d N_OUT7_Mp8@94_g N_VDD_Mp8@94_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@93 N_OUT8_Mn8@93_d N_OUT7_Mn8@93_g N_VSS_Mn8@93_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@92 N_OUT8_Mn8@92_d N_OUT7_Mn8@92_g N_VSS_Mn8@92_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@93 N_OUT8_Mp8@93_d N_OUT7_Mp8@93_g N_VDD_Mp8@93_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@92 N_OUT8_Mp8@92_d N_OUT7_Mp8@92_g N_VDD_Mp8@92_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@91 N_OUT8_Mn8@91_d N_OUT7_Mn8@91_g N_VSS_Mn8@91_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@90 N_OUT8_Mn8@90_d N_OUT7_Mn8@90_g N_VSS_Mn8@90_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@91 N_OUT8_Mp8@91_d N_OUT7_Mp8@91_g N_VDD_Mp8@91_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@90 N_OUT8_Mp8@90_d N_OUT7_Mp8@90_g N_VDD_Mp8@90_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@89 N_OUT8_Mn8@89_d N_OUT7_Mn8@89_g N_VSS_Mn8@89_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@88 N_OUT8_Mn8@88_d N_OUT7_Mn8@88_g N_VSS_Mn8@88_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@89 N_OUT8_Mp8@89_d N_OUT7_Mp8@89_g N_VDD_Mp8@89_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@88 N_OUT8_Mp8@88_d N_OUT7_Mp8@88_g N_VDD_Mp8@88_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@87 N_OUT8_Mn8@87_d N_OUT7_Mn8@87_g N_VSS_Mn8@87_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@86 N_OUT8_Mn8@86_d N_OUT7_Mn8@86_g N_VSS_Mn8@86_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@87 N_OUT8_Mp8@87_d N_OUT7_Mp8@87_g N_VDD_Mp8@87_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@86 N_OUT8_Mp8@86_d N_OUT7_Mp8@86_g N_VDD_Mp8@86_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@85 N_OUT8_Mn8@85_d N_OUT7_Mn8@85_g N_VSS_Mn8@85_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@84 N_OUT8_Mn8@84_d N_OUT7_Mn8@84_g N_VSS_Mn8@84_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@85 N_OUT8_Mp8@85_d N_OUT7_Mp8@85_g N_VDD_Mp8@85_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@84 N_OUT8_Mp8@84_d N_OUT7_Mp8@84_g N_VDD_Mp8@84_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@83 N_OUT8_Mn8@83_d N_OUT7_Mn8@83_g N_VSS_Mn8@83_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@82 N_OUT8_Mn8@82_d N_OUT7_Mn8@82_g N_VSS_Mn8@82_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@83 N_OUT8_Mp8@83_d N_OUT7_Mp8@83_g N_VDD_Mp8@83_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@82 N_OUT8_Mp8@82_d N_OUT7_Mp8@82_g N_VDD_Mp8@82_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@81 N_OUT8_Mn8@81_d N_OUT7_Mn8@81_g N_VSS_Mn8@81_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@80 N_OUT8_Mn8@80_d N_OUT7_Mn8@80_g N_VSS_Mn8@80_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@81 N_OUT8_Mp8@81_d N_OUT7_Mp8@81_g N_VDD_Mp8@81_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@80 N_OUT8_Mp8@80_d N_OUT7_Mp8@80_g N_VDD_Mp8@80_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@79 N_OUT8_Mn8@79_d N_OUT7_Mn8@79_g N_VSS_Mn8@79_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@78 N_OUT8_Mn8@78_d N_OUT7_Mn8@78_g N_VSS_Mn8@78_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@79 N_OUT8_Mp8@79_d N_OUT7_Mp8@79_g N_VDD_Mp8@79_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@78 N_OUT8_Mp8@78_d N_OUT7_Mp8@78_g N_VDD_Mp8@78_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@77 N_OUT8_Mn8@77_d N_OUT7_Mn8@77_g N_VSS_Mn8@77_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@76 N_OUT8_Mn8@76_d N_OUT7_Mn8@76_g N_VSS_Mn8@76_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@77 N_OUT8_Mp8@77_d N_OUT7_Mp8@77_g N_VDD_Mp8@77_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@76 N_OUT8_Mp8@76_d N_OUT7_Mp8@76_g N_VDD_Mp8@76_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@75 N_OUT8_Mn8@75_d N_OUT7_Mn8@75_g N_VSS_Mn8@75_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@74 N_OUT8_Mn8@74_d N_OUT7_Mn8@74_g N_VSS_Mn8@74_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@75 N_OUT8_Mp8@75_d N_OUT7_Mp8@75_g N_VDD_Mp8@75_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@74 N_OUT8_Mp8@74_d N_OUT7_Mp8@74_g N_VDD_Mp8@74_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@73 N_OUT8_Mn8@73_d N_OUT7_Mn8@73_g N_VSS_Mn8@73_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@72 N_OUT8_Mn8@72_d N_OUT7_Mn8@72_g N_VSS_Mn8@72_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@73 N_OUT8_Mp8@73_d N_OUT7_Mp8@73_g N_VDD_Mp8@73_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@72 N_OUT8_Mp8@72_d N_OUT7_Mp8@72_g N_VDD_Mp8@72_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@71 N_OUT8_Mn8@71_d N_OUT7_Mn8@71_g N_VSS_Mn8@71_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@70 N_OUT8_Mn8@70_d N_OUT7_Mn8@70_g N_VSS_Mn8@70_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@71 N_OUT8_Mp8@71_d N_OUT7_Mp8@71_g N_VDD_Mp8@71_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@70 N_OUT8_Mp8@70_d N_OUT7_Mp8@70_g N_VDD_Mp8@70_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@69 N_OUT8_Mn8@69_d N_OUT7_Mn8@69_g N_VSS_Mn8@69_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@68 N_OUT8_Mn8@68_d N_OUT7_Mn8@68_g N_VSS_Mn8@68_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@69 N_OUT8_Mp8@69_d N_OUT7_Mp8@69_g N_VDD_Mp8@69_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@68 N_OUT8_Mp8@68_d N_OUT7_Mp8@68_g N_VDD_Mp8@68_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@67 N_OUT8_Mn8@67_d N_OUT7_Mn8@67_g N_VSS_Mn8@67_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@66 N_OUT8_Mn8@66_d N_OUT7_Mn8@66_g N_VSS_Mn8@66_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@67 N_OUT8_Mp8@67_d N_OUT7_Mp8@67_g N_VDD_Mp8@67_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@66 N_OUT8_Mp8@66_d N_OUT7_Mp8@66_g N_VDD_Mp8@66_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@65 N_OUT8_Mn8@65_d N_OUT7_Mn8@65_g N_VSS_Mn8@65_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@64 N_OUT8_Mn8@64_d N_OUT7_Mn8@64_g N_VSS_Mn8@64_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@65 N_OUT8_Mp8@65_d N_OUT7_Mp8@65_g N_VDD_Mp8@65_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@64 N_OUT8_Mp8@64_d N_OUT7_Mp8@64_g N_VDD_Mp8@64_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@63 N_OUT8_Mn8@63_d N_OUT7_Mn8@63_g N_VSS_Mn8@63_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@62 N_OUT8_Mn8@62_d N_OUT7_Mn8@62_g N_VSS_Mn8@62_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@63 N_OUT8_Mp8@63_d N_OUT7_Mp8@63_g N_VDD_Mp8@63_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@62 N_OUT8_Mp8@62_d N_OUT7_Mp8@62_g N_VDD_Mp8@62_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@61 N_OUT8_Mn8@61_d N_OUT7_Mn8@61_g N_VSS_Mn8@61_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@60 N_OUT8_Mn8@60_d N_OUT7_Mn8@60_g N_VSS_Mn8@60_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@61 N_OUT8_Mp8@61_d N_OUT7_Mp8@61_g N_VDD_Mp8@61_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@60 N_OUT8_Mp8@60_d N_OUT7_Mp8@60_g N_VDD_Mp8@60_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@59 N_OUT8_Mn8@59_d N_OUT7_Mn8@59_g N_VSS_Mn8@59_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@58 N_OUT8_Mn8@58_d N_OUT7_Mn8@58_g N_VSS_Mn8@58_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@59 N_OUT8_Mp8@59_d N_OUT7_Mp8@59_g N_VDD_Mp8@59_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@58 N_OUT8_Mp8@58_d N_OUT7_Mp8@58_g N_VDD_Mp8@58_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@57 N_OUT8_Mn8@57_d N_OUT7_Mn8@57_g N_VSS_Mn8@57_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@56 N_OUT8_Mn8@56_d N_OUT7_Mn8@56_g N_VSS_Mn8@56_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@57 N_OUT8_Mp8@57_d N_OUT7_Mp8@57_g N_VDD_Mp8@57_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@56 N_OUT8_Mp8@56_d N_OUT7_Mp8@56_g N_VDD_Mp8@56_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@55 N_OUT8_Mn8@55_d N_OUT7_Mn8@55_g N_VSS_Mn8@55_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@54 N_OUT8_Mn8@54_d N_OUT7_Mn8@54_g N_VSS_Mn8@54_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@55 N_OUT8_Mp8@55_d N_OUT7_Mp8@55_g N_VDD_Mp8@55_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@54 N_OUT8_Mp8@54_d N_OUT7_Mp8@54_g N_VDD_Mp8@54_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@53 N_OUT8_Mn8@53_d N_OUT7_Mn8@53_g N_VSS_Mn8@53_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@52 N_OUT8_Mn8@52_d N_OUT7_Mn8@52_g N_VSS_Mn8@52_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@53 N_OUT8_Mp8@53_d N_OUT7_Mp8@53_g N_VDD_Mp8@53_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@52 N_OUT8_Mp8@52_d N_OUT7_Mp8@52_g N_VDD_Mp8@52_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@51 N_OUT8_Mn8@51_d N_OUT7_Mn8@51_g N_VSS_Mn8@51_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@50 N_OUT8_Mn8@50_d N_OUT7_Mn8@50_g N_VSS_Mn8@50_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@51 N_OUT8_Mp8@51_d N_OUT7_Mp8@51_g N_VDD_Mp8@51_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@50 N_OUT8_Mp8@50_d N_OUT7_Mp8@50_g N_VDD_Mp8@50_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@49 N_OUT8_Mn8@49_d N_OUT7_Mn8@49_g N_VSS_Mn8@49_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@48 N_OUT8_Mn8@48_d N_OUT7_Mn8@48_g N_VSS_Mn8@48_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@49 N_OUT8_Mp8@49_d N_OUT7_Mp8@49_g N_VDD_Mp8@49_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@48 N_OUT8_Mp8@48_d N_OUT7_Mp8@48_g N_VDD_Mp8@48_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@47 N_OUT8_Mn8@47_d N_OUT7_Mn8@47_g N_VSS_Mn8@47_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@46 N_OUT8_Mn8@46_d N_OUT7_Mn8@46_g N_VSS_Mn8@46_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@47 N_OUT8_Mp8@47_d N_OUT7_Mp8@47_g N_VDD_Mp8@47_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@46 N_OUT8_Mp8@46_d N_OUT7_Mp8@46_g N_VDD_Mp8@46_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@45 N_OUT8_Mn8@45_d N_OUT7_Mn8@45_g N_VSS_Mn8@45_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@44 N_OUT8_Mn8@44_d N_OUT7_Mn8@44_g N_VSS_Mn8@44_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@45 N_OUT8_Mp8@45_d N_OUT7_Mp8@45_g N_VDD_Mp8@45_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@44 N_OUT8_Mp8@44_d N_OUT7_Mp8@44_g N_VDD_Mp8@44_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@43 N_OUT8_Mn8@43_d N_OUT7_Mn8@43_g N_VSS_Mn8@43_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@42 N_OUT8_Mn8@42_d N_OUT7_Mn8@42_g N_VSS_Mn8@42_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@43 N_OUT8_Mp8@43_d N_OUT7_Mp8@43_g N_VDD_Mp8@43_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@42 N_OUT8_Mp8@42_d N_OUT7_Mp8@42_g N_VDD_Mp8@42_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@41 N_OUT8_Mn8@41_d N_OUT7_Mn8@41_g N_VSS_Mn8@41_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@40 N_OUT8_Mn8@40_d N_OUT7_Mn8@40_g N_VSS_Mn8@40_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@41 N_OUT8_Mp8@41_d N_OUT7_Mp8@41_g N_VDD_Mp8@41_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@40 N_OUT8_Mp8@40_d N_OUT7_Mp8@40_g N_VDD_Mp8@40_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@39 N_OUT8_Mn8@39_d N_OUT7_Mn8@39_g N_VSS_Mn8@39_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@38 N_OUT8_Mn8@38_d N_OUT7_Mn8@38_g N_VSS_Mn8@38_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@39 N_OUT8_Mp8@39_d N_OUT7_Mp8@39_g N_VDD_Mp8@39_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@38 N_OUT8_Mp8@38_d N_OUT7_Mp8@38_g N_VDD_Mp8@38_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@37 N_OUT8_Mn8@37_d N_OUT7_Mn8@37_g N_VSS_Mn8@37_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@36 N_OUT8_Mn8@36_d N_OUT7_Mn8@36_g N_VSS_Mn8@36_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@37 N_OUT8_Mp8@37_d N_OUT7_Mp8@37_g N_VDD_Mp8@37_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@36 N_OUT8_Mp8@36_d N_OUT7_Mp8@36_g N_VDD_Mp8@36_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@35 N_OUT8_Mn8@35_d N_OUT7_Mn8@35_g N_VSS_Mn8@35_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@34 N_OUT8_Mn8@34_d N_OUT7_Mn8@34_g N_VSS_Mn8@34_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@35 N_OUT8_Mp8@35_d N_OUT7_Mp8@35_g N_VDD_Mp8@35_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@34 N_OUT8_Mp8@34_d N_OUT7_Mp8@34_g N_VDD_Mp8@34_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@33 N_OUT8_Mn8@33_d N_OUT7_Mn8@33_g N_VSS_Mn8@33_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@32 N_OUT8_Mn8@32_d N_OUT7_Mn8@32_g N_VSS_Mn8@32_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@33 N_OUT8_Mp8@33_d N_OUT7_Mp8@33_g N_VDD_Mp8@33_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@32 N_OUT8_Mp8@32_d N_OUT7_Mp8@32_g N_VDD_Mp8@32_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@31 N_OUT8_Mn8@31_d N_OUT7_Mn8@31_g N_VSS_Mn8@31_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@30 N_OUT8_Mn8@30_d N_OUT7_Mn8@30_g N_VSS_Mn8@30_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@31 N_OUT8_Mp8@31_d N_OUT7_Mp8@31_g N_VDD_Mp8@31_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@30 N_OUT8_Mp8@30_d N_OUT7_Mp8@30_g N_VDD_Mp8@30_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@29 N_OUT8_Mn8@29_d N_OUT7_Mn8@29_g N_VSS_Mn8@29_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@28 N_OUT8_Mn8@28_d N_OUT7_Mn8@28_g N_VSS_Mn8@28_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@29 N_OUT8_Mp8@29_d N_OUT7_Mp8@29_g N_VDD_Mp8@29_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@28 N_OUT8_Mp8@28_d N_OUT7_Mp8@28_g N_VDD_Mp8@28_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@27 N_OUT8_Mn8@27_d N_OUT7_Mn8@27_g N_VSS_Mn8@27_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@26 N_OUT8_Mn8@26_d N_OUT7_Mn8@26_g N_VSS_Mn8@26_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@27 N_OUT8_Mp8@27_d N_OUT7_Mp8@27_g N_VDD_Mp8@27_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@26 N_OUT8_Mp8@26_d N_OUT7_Mp8@26_g N_VDD_Mp8@26_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@25 N_OUT8_Mn8@25_d N_OUT7_Mn8@25_g N_VSS_Mn8@25_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@24 N_OUT8_Mn8@24_d N_OUT7_Mn8@24_g N_VSS_Mn8@24_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@25 N_OUT8_Mp8@25_d N_OUT7_Mp8@25_g N_VDD_Mp8@25_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@24 N_OUT8_Mp8@24_d N_OUT7_Mp8@24_g N_VDD_Mp8@24_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@23 N_OUT8_Mn8@23_d N_OUT7_Mn8@23_g N_VSS_Mn8@23_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@22 N_OUT8_Mn8@22_d N_OUT7_Mn8@22_g N_VSS_Mn8@22_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@23 N_OUT8_Mp8@23_d N_OUT7_Mp8@23_g N_VDD_Mp8@23_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@22 N_OUT8_Mp8@22_d N_OUT7_Mp8@22_g N_VDD_Mp8@22_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@21 N_OUT8_Mn8@21_d N_OUT7_Mn8@21_g N_VSS_Mn8@21_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@20 N_OUT8_Mn8@20_d N_OUT7_Mn8@20_g N_VSS_Mn8@20_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@21 N_OUT8_Mp8@21_d N_OUT7_Mp8@21_g N_VDD_Mp8@21_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@20 N_OUT8_Mp8@20_d N_OUT7_Mp8@20_g N_VDD_Mp8@20_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@19 N_OUT8_Mn8@19_d N_OUT7_Mn8@19_g N_VSS_Mn8@19_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@18 N_OUT8_Mn8@18_d N_OUT7_Mn8@18_g N_VSS_Mn8@18_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@19 N_OUT8_Mp8@19_d N_OUT7_Mp8@19_g N_VDD_Mp8@19_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@18 N_OUT8_Mp8@18_d N_OUT7_Mp8@18_g N_VDD_Mp8@18_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@17 N_OUT8_Mn8@17_d N_OUT7_Mn8@17_g N_VSS_Mn8@17_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@16 N_OUT8_Mn8@16_d N_OUT7_Mn8@16_g N_VSS_Mn8@16_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@17 N_OUT8_Mp8@17_d N_OUT7_Mp8@17_g N_VDD_Mp8@17_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@16 N_OUT8_Mp8@16_d N_OUT7_Mp8@16_g N_VDD_Mp8@16_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@15 N_OUT8_Mn8@15_d N_OUT7_Mn8@15_g N_VSS_Mn8@15_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@14 N_OUT8_Mn8@14_d N_OUT7_Mn8@14_g N_VSS_Mn8@14_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@15 N_OUT8_Mp8@15_d N_OUT7_Mp8@15_g N_VDD_Mp8@15_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@14 N_OUT8_Mp8@14_d N_OUT7_Mp8@14_g N_VDD_Mp8@14_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@13 N_OUT8_Mn8@13_d N_OUT7_Mn8@13_g N_VSS_Mn8@13_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@12 N_OUT8_Mn8@12_d N_OUT7_Mn8@12_g N_VSS_Mn8@12_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@13 N_OUT8_Mp8@13_d N_OUT7_Mp8@13_g N_VDD_Mp8@13_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@12 N_OUT8_Mp8@12_d N_OUT7_Mp8@12_g N_VDD_Mp8@12_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@11 N_OUT8_Mn8@11_d N_OUT7_Mn8@11_g N_VSS_Mn8@11_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@10 N_OUT8_Mn8@10_d N_OUT7_Mn8@10_g N_VSS_Mn8@10_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@11 N_OUT8_Mp8@11_d N_OUT7_Mp8@11_g N_VDD_Mp8@11_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@10 N_OUT8_Mp8@10_d N_OUT7_Mp8@10_g N_VDD_Mp8@10_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@9 N_OUT8_Mn8@9_d N_OUT7_Mn8@9_g N_VSS_Mn8@9_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@8 N_OUT8_Mn8@8_d N_OUT7_Mn8@8_g N_VSS_Mn8@8_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@9 N_OUT8_Mp8@9_d N_OUT7_Mp8@9_g N_VDD_Mp8@9_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@8 N_OUT8_Mp8@8_d N_OUT7_Mp8@8_g N_VDD_Mp8@8_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@7 N_OUT8_Mn8@7_d N_OUT7_Mn8@7_g N_VSS_Mn8@7_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@6 N_OUT8_Mn8@6_d N_OUT7_Mn8@6_g N_VSS_Mn8@6_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@7 N_OUT8_Mp8@7_d N_OUT7_Mp8@7_g N_VDD_Mp8@7_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@6 N_OUT8_Mp8@6_d N_OUT7_Mp8@6_g N_VDD_Mp8@6_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@5 N_OUT8_Mn8@5_d N_OUT7_Mn8@5_g N_VSS_Mn8@5_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@4 N_OUT8_Mn8@4_d N_OUT7_Mn8@4_g N_VSS_Mn8@4_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@5 N_OUT8_Mp8@5_d N_OUT7_Mp8@5_g N_VDD_Mp8@5_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@4 N_OUT8_Mp8@4_d N_OUT7_Mp8@4_g N_VDD_Mp8@4_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn8@3 N_OUT8_Mn8@3_d N_OUT7_Mn8@3_g N_VSS_Mn8@3_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mn8@2 N_OUT8_Mn8@2_d N_OUT7_Mn8@2_g N_VSS_Mn8@2_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=5e-07 AD=1.325e-13 AS=1.4125e-13 PD=5.3e-07 PS=5.65e-07
Mp8@3 N_OUT8_Mp8@3_d N_OUT7_Mp8@3_g N_VDD_Mp8@3_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mp8@2 N_OUT8_Mp8@2_d N_OUT7_Mp8@2_g N_VDD_Mp8@2_s N_VDD_Mp8@3769_b P_18
+ L=1.8e-07 W=1.5e-06 AD=3.9375e-13 AS=4.275e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4097 N_OUT9_Mn9@4097_d N_OUT8_Mn9@4097_g N_VSS_Mn9@4097_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4096 N_OUT9_Mn9@4096_d N_OUT8_Mn9@4096_g N_VSS_Mn9@4096_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4097 N_OUT9_Mp9@4097_d N_OUT8_Mp9@4097_g N_VDD_Mp9@4097_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4096 N_OUT9_Mp9@4096_d N_OUT8_Mp9@4096_g N_VDD_Mp9@4096_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4095 N_OUT9_Mn9@4095_d N_OUT8_Mn9@4095_g N_VSS_Mn9@4095_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4094 N_OUT9_Mn9@4094_d N_OUT8_Mn9@4094_g N_VSS_Mn9@4094_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4095 N_OUT9_Mp9@4095_d N_OUT8_Mp9@4095_g N_VDD_Mp9@4095_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4094 N_OUT9_Mp9@4094_d N_OUT8_Mp9@4094_g N_VDD_Mp9@4094_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4093 N_OUT9_Mn9@4093_d N_OUT8_Mn9@4093_g N_VSS_Mn9@4093_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4092 N_OUT9_Mn9@4092_d N_OUT8_Mn9@4092_g N_VSS_Mn9@4092_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4093 N_OUT9_Mp9@4093_d N_OUT8_Mp9@4093_g N_VDD_Mp9@4093_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4092 N_OUT9_Mp9@4092_d N_OUT8_Mp9@4092_g N_VDD_Mp9@4092_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4091 N_OUT9_Mn9@4091_d N_OUT8_Mn9@4091_g N_VSS_Mn9@4091_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4090 N_OUT9_Mn9@4090_d N_OUT8_Mn9@4090_g N_VSS_Mn9@4090_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4091 N_OUT9_Mp9@4091_d N_OUT8_Mp9@4091_g N_VDD_Mp9@4091_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4090 N_OUT9_Mp9@4090_d N_OUT8_Mp9@4090_g N_VDD_Mp9@4090_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4089 N_OUT9_Mn9@4089_d N_OUT8_Mn9@4089_g N_VSS_Mn9@4089_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4088 N_OUT9_Mn9@4088_d N_OUT8_Mn9@4088_g N_VSS_Mn9@4088_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4089 N_OUT9_Mp9@4089_d N_OUT8_Mp9@4089_g N_VDD_Mp9@4089_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4088 N_OUT9_Mp9@4088_d N_OUT8_Mp9@4088_g N_VDD_Mp9@4088_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4087 N_OUT9_Mn9@4087_d N_OUT8_Mn9@4087_g N_VSS_Mn9@4087_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4086 N_OUT9_Mn9@4086_d N_OUT8_Mn9@4086_g N_VSS_Mn9@4086_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4087 N_OUT9_Mp9@4087_d N_OUT8_Mp9@4087_g N_VDD_Mp9@4087_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4086 N_OUT9_Mp9@4086_d N_OUT8_Mp9@4086_g N_VDD_Mp9@4086_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4085 N_OUT9_Mn9@4085_d N_OUT8_Mn9@4085_g N_VSS_Mn9@4085_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4084 N_OUT9_Mn9@4084_d N_OUT8_Mn9@4084_g N_VSS_Mn9@4084_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4085 N_OUT9_Mp9@4085_d N_OUT8_Mp9@4085_g N_VDD_Mp9@4085_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4084 N_OUT9_Mp9@4084_d N_OUT8_Mp9@4084_g N_VDD_Mp9@4084_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4083 N_OUT9_Mn9@4083_d N_OUT8_Mn9@4083_g N_VSS_Mn9@4083_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4082 N_OUT9_Mn9@4082_d N_OUT8_Mn9@4082_g N_VSS_Mn9@4082_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4083 N_OUT9_Mp9@4083_d N_OUT8_Mp9@4083_g N_VDD_Mp9@4083_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4082 N_OUT9_Mp9@4082_d N_OUT8_Mp9@4082_g N_VDD_Mp9@4082_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4081 N_OUT9_Mn9@4081_d N_OUT8_Mn9@4081_g N_VSS_Mn9@4081_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4080 N_OUT9_Mn9@4080_d N_OUT8_Mn9@4080_g N_VSS_Mn9@4080_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4081 N_OUT9_Mp9@4081_d N_OUT8_Mp9@4081_g N_VDD_Mp9@4081_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4080 N_OUT9_Mp9@4080_d N_OUT8_Mp9@4080_g N_VDD_Mp9@4080_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4079 N_OUT9_Mn9@4079_d N_OUT8_Mn9@4079_g N_VSS_Mn9@4079_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4078 N_OUT9_Mn9@4078_d N_OUT8_Mn9@4078_g N_VSS_Mn9@4078_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4079 N_OUT9_Mp9@4079_d N_OUT8_Mp9@4079_g N_VDD_Mp9@4079_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4078 N_OUT9_Mp9@4078_d N_OUT8_Mp9@4078_g N_VDD_Mp9@4078_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4077 N_OUT9_Mn9@4077_d N_OUT8_Mn9@4077_g N_VSS_Mn9@4077_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4076 N_OUT9_Mn9@4076_d N_OUT8_Mn9@4076_g N_VSS_Mn9@4076_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4077 N_OUT9_Mp9@4077_d N_OUT8_Mp9@4077_g N_VDD_Mp9@4077_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4076 N_OUT9_Mp9@4076_d N_OUT8_Mp9@4076_g N_VDD_Mp9@4076_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4075 N_OUT9_Mn9@4075_d N_OUT8_Mn9@4075_g N_VSS_Mn9@4075_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4074 N_OUT9_Mn9@4074_d N_OUT8_Mn9@4074_g N_VSS_Mn9@4074_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4075 N_OUT9_Mp9@4075_d N_OUT8_Mp9@4075_g N_VDD_Mp9@4075_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4074 N_OUT9_Mp9@4074_d N_OUT8_Mp9@4074_g N_VDD_Mp9@4074_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4073 N_OUT9_Mn9@4073_d N_OUT8_Mn9@4073_g N_VSS_Mn9@4073_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4072 N_OUT9_Mn9@4072_d N_OUT8_Mn9@4072_g N_VSS_Mn9@4072_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4073 N_OUT9_Mp9@4073_d N_OUT8_Mp9@4073_g N_VDD_Mp9@4073_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4072 N_OUT9_Mp9@4072_d N_OUT8_Mp9@4072_g N_VDD_Mp9@4072_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4071 N_OUT9_Mn9@4071_d N_OUT8_Mn9@4071_g N_VSS_Mn9@4071_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4070 N_OUT9_Mn9@4070_d N_OUT8_Mn9@4070_g N_VSS_Mn9@4070_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4071 N_OUT9_Mp9@4071_d N_OUT8_Mp9@4071_g N_VDD_Mp9@4071_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4070 N_OUT9_Mp9@4070_d N_OUT8_Mp9@4070_g N_VDD_Mp9@4070_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4069 N_OUT9_Mn9@4069_d N_OUT8_Mn9@4069_g N_VSS_Mn9@4069_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4068 N_OUT9_Mn9@4068_d N_OUT8_Mn9@4068_g N_VSS_Mn9@4068_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4069 N_OUT9_Mp9@4069_d N_OUT8_Mp9@4069_g N_VDD_Mp9@4069_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4068 N_OUT9_Mp9@4068_d N_OUT8_Mp9@4068_g N_VDD_Mp9@4068_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4067 N_OUT9_Mn9@4067_d N_OUT8_Mn9@4067_g N_VSS_Mn9@4067_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4066 N_OUT9_Mn9@4066_d N_OUT8_Mn9@4066_g N_VSS_Mn9@4066_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4067 N_OUT9_Mp9@4067_d N_OUT8_Mp9@4067_g N_VDD_Mp9@4067_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4066 N_OUT9_Mp9@4066_d N_OUT8_Mp9@4066_g N_VDD_Mp9@4066_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4065 N_OUT9_Mn9@4065_d N_OUT8_Mn9@4065_g N_VSS_Mn9@4065_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4064 N_OUT9_Mn9@4064_d N_OUT8_Mn9@4064_g N_VSS_Mn9@4064_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4065 N_OUT9_Mp9@4065_d N_OUT8_Mp9@4065_g N_VDD_Mp9@4065_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4064 N_OUT9_Mp9@4064_d N_OUT8_Mp9@4064_g N_VDD_Mp9@4064_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4063 N_OUT9_Mn9@4063_d N_OUT8_Mn9@4063_g N_VSS_Mn9@4063_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4062 N_OUT9_Mn9@4062_d N_OUT8_Mn9@4062_g N_VSS_Mn9@4062_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4063 N_OUT9_Mp9@4063_d N_OUT8_Mp9@4063_g N_VDD_Mp9@4063_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4062 N_OUT9_Mp9@4062_d N_OUT8_Mp9@4062_g N_VDD_Mp9@4062_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4061 N_OUT9_Mn9@4061_d N_OUT8_Mn9@4061_g N_VSS_Mn9@4061_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4060 N_OUT9_Mn9@4060_d N_OUT8_Mn9@4060_g N_VSS_Mn9@4060_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4061 N_OUT9_Mp9@4061_d N_OUT8_Mp9@4061_g N_VDD_Mp9@4061_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4060 N_OUT9_Mp9@4060_d N_OUT8_Mp9@4060_g N_VDD_Mp9@4060_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4059 N_OUT9_Mn9@4059_d N_OUT8_Mn9@4059_g N_VSS_Mn9@4059_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4058 N_OUT9_Mn9@4058_d N_OUT8_Mn9@4058_g N_VSS_Mn9@4058_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4059 N_OUT9_Mp9@4059_d N_OUT8_Mp9@4059_g N_VDD_Mp9@4059_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4058 N_OUT9_Mp9@4058_d N_OUT8_Mp9@4058_g N_VDD_Mp9@4058_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4057 N_OUT9_Mn9@4057_d N_OUT8_Mn9@4057_g N_VSS_Mn9@4057_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4056 N_OUT9_Mn9@4056_d N_OUT8_Mn9@4056_g N_VSS_Mn9@4056_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4057 N_OUT9_Mp9@4057_d N_OUT8_Mp9@4057_g N_VDD_Mp9@4057_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4056 N_OUT9_Mp9@4056_d N_OUT8_Mp9@4056_g N_VDD_Mp9@4056_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4055 N_OUT9_Mn9@4055_d N_OUT8_Mn9@4055_g N_VSS_Mn9@4055_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4054 N_OUT9_Mn9@4054_d N_OUT8_Mn9@4054_g N_VSS_Mn9@4054_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4055 N_OUT9_Mp9@4055_d N_OUT8_Mp9@4055_g N_VDD_Mp9@4055_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4054 N_OUT9_Mp9@4054_d N_OUT8_Mp9@4054_g N_VDD_Mp9@4054_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4053 N_OUT9_Mn9@4053_d N_OUT8_Mn9@4053_g N_VSS_Mn9@4053_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4052 N_OUT9_Mn9@4052_d N_OUT8_Mn9@4052_g N_VSS_Mn9@4052_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4053 N_OUT9_Mp9@4053_d N_OUT8_Mp9@4053_g N_VDD_Mp9@4053_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4052 N_OUT9_Mp9@4052_d N_OUT8_Mp9@4052_g N_VDD_Mp9@4052_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4051 N_OUT9_Mn9@4051_d N_OUT8_Mn9@4051_g N_VSS_Mn9@4051_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4050 N_OUT9_Mn9@4050_d N_OUT8_Mn9@4050_g N_VSS_Mn9@4050_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4051 N_OUT9_Mp9@4051_d N_OUT8_Mp9@4051_g N_VDD_Mp9@4051_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4050 N_OUT9_Mp9@4050_d N_OUT8_Mp9@4050_g N_VDD_Mp9@4050_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4049 N_OUT9_Mn9@4049_d N_OUT8_Mn9@4049_g N_VSS_Mn9@4049_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4048 N_OUT9_Mn9@4048_d N_OUT8_Mn9@4048_g N_VSS_Mn9@4048_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4049 N_OUT9_Mp9@4049_d N_OUT8_Mp9@4049_g N_VDD_Mp9@4049_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4048 N_OUT9_Mp9@4048_d N_OUT8_Mp9@4048_g N_VDD_Mp9@4048_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4047 N_OUT9_Mn9@4047_d N_OUT8_Mn9@4047_g N_VSS_Mn9@4047_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4046 N_OUT9_Mn9@4046_d N_OUT8_Mn9@4046_g N_VSS_Mn9@4046_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4047 N_OUT9_Mp9@4047_d N_OUT8_Mp9@4047_g N_VDD_Mp9@4047_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4046 N_OUT9_Mp9@4046_d N_OUT8_Mp9@4046_g N_VDD_Mp9@4046_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4045 N_OUT9_Mn9@4045_d N_OUT8_Mn9@4045_g N_VSS_Mn9@4045_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4044 N_OUT9_Mn9@4044_d N_OUT8_Mn9@4044_g N_VSS_Mn9@4044_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4045 N_OUT9_Mp9@4045_d N_OUT8_Mp9@4045_g N_VDD_Mp9@4045_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4044 N_OUT9_Mp9@4044_d N_OUT8_Mp9@4044_g N_VDD_Mp9@4044_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4043 N_OUT9_Mn9@4043_d N_OUT8_Mn9@4043_g N_VSS_Mn9@4043_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4042 N_OUT9_Mn9@4042_d N_OUT8_Mn9@4042_g N_VSS_Mn9@4042_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4043 N_OUT9_Mp9@4043_d N_OUT8_Mp9@4043_g N_VDD_Mp9@4043_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4042 N_OUT9_Mp9@4042_d N_OUT8_Mp9@4042_g N_VDD_Mp9@4042_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4041 N_OUT9_Mn9@4041_d N_OUT8_Mn9@4041_g N_VSS_Mn9@4041_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4040 N_OUT9_Mn9@4040_d N_OUT8_Mn9@4040_g N_VSS_Mn9@4040_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4041 N_OUT9_Mp9@4041_d N_OUT8_Mp9@4041_g N_VDD_Mp9@4041_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4040 N_OUT9_Mp9@4040_d N_OUT8_Mp9@4040_g N_VDD_Mp9@4040_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4039 N_OUT9_Mn9@4039_d N_OUT8_Mn9@4039_g N_VSS_Mn9@4039_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4038 N_OUT9_Mn9@4038_d N_OUT8_Mn9@4038_g N_VSS_Mn9@4038_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4039 N_OUT9_Mp9@4039_d N_OUT8_Mp9@4039_g N_VDD_Mp9@4039_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4038 N_OUT9_Mp9@4038_d N_OUT8_Mp9@4038_g N_VDD_Mp9@4038_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4037 N_OUT9_Mn9@4037_d N_OUT8_Mn9@4037_g N_VSS_Mn9@4037_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4036 N_OUT9_Mn9@4036_d N_OUT8_Mn9@4036_g N_VSS_Mn9@4036_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4037 N_OUT9_Mp9@4037_d N_OUT8_Mp9@4037_g N_VDD_Mp9@4037_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4036 N_OUT9_Mp9@4036_d N_OUT8_Mp9@4036_g N_VDD_Mp9@4036_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4035 N_OUT9_Mn9@4035_d N_OUT8_Mn9@4035_g N_VSS_Mn9@4035_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4034 N_OUT9_Mn9@4034_d N_OUT8_Mn9@4034_g N_VSS_Mn9@4034_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4035 N_OUT9_Mp9@4035_d N_OUT8_Mp9@4035_g N_VDD_Mp9@4035_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4034 N_OUT9_Mp9@4034_d N_OUT8_Mp9@4034_g N_VDD_Mp9@4034_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4033 N_OUT9_Mn9@4033_d N_OUT8_Mn9@4033_g N_VSS_Mn9@4033_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4032 N_OUT9_Mn9@4032_d N_OUT8_Mn9@4032_g N_VSS_Mn9@4032_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4033 N_OUT9_Mp9@4033_d N_OUT8_Mp9@4033_g N_VDD_Mp9@4033_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4032 N_OUT9_Mp9@4032_d N_OUT8_Mp9@4032_g N_VDD_Mp9@4032_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4031 N_OUT9_Mn9@4031_d N_OUT8_Mn9@4031_g N_VSS_Mn9@4031_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4030 N_OUT9_Mn9@4030_d N_OUT8_Mn9@4030_g N_VSS_Mn9@4030_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4031 N_OUT9_Mp9@4031_d N_OUT8_Mp9@4031_g N_VDD_Mp9@4031_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4030 N_OUT9_Mp9@4030_d N_OUT8_Mp9@4030_g N_VDD_Mp9@4030_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4029 N_OUT9_Mn9@4029_d N_OUT8_Mn9@4029_g N_VSS_Mn9@4029_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4028 N_OUT9_Mn9@4028_d N_OUT8_Mn9@4028_g N_VSS_Mn9@4028_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4029 N_OUT9_Mp9@4029_d N_OUT8_Mp9@4029_g N_VDD_Mp9@4029_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4028 N_OUT9_Mp9@4028_d N_OUT8_Mp9@4028_g N_VDD_Mp9@4028_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4027 N_OUT9_Mn9@4027_d N_OUT8_Mn9@4027_g N_VSS_Mn9@4027_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4026 N_OUT9_Mn9@4026_d N_OUT8_Mn9@4026_g N_VSS_Mn9@4026_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4027 N_OUT9_Mp9@4027_d N_OUT8_Mp9@4027_g N_VDD_Mp9@4027_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4026 N_OUT9_Mp9@4026_d N_OUT8_Mp9@4026_g N_VDD_Mp9@4026_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4025 N_OUT9_Mn9@4025_d N_OUT8_Mn9@4025_g N_VSS_Mn9@4025_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4024 N_OUT9_Mn9@4024_d N_OUT8_Mn9@4024_g N_VSS_Mn9@4024_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4025 N_OUT9_Mp9@4025_d N_OUT8_Mp9@4025_g N_VDD_Mp9@4025_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4024 N_OUT9_Mp9@4024_d N_OUT8_Mp9@4024_g N_VDD_Mp9@4024_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4023 N_OUT9_Mn9@4023_d N_OUT8_Mn9@4023_g N_VSS_Mn9@4023_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4022 N_OUT9_Mn9@4022_d N_OUT8_Mn9@4022_g N_VSS_Mn9@4022_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4023 N_OUT9_Mp9@4023_d N_OUT8_Mp9@4023_g N_VDD_Mp9@4023_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4022 N_OUT9_Mp9@4022_d N_OUT8_Mp9@4022_g N_VDD_Mp9@4022_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4021 N_OUT9_Mn9@4021_d N_OUT8_Mn9@4021_g N_VSS_Mn9@4021_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4020 N_OUT9_Mn9@4020_d N_OUT8_Mn9@4020_g N_VSS_Mn9@4020_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4021 N_OUT9_Mp9@4021_d N_OUT8_Mp9@4021_g N_VDD_Mp9@4021_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4020 N_OUT9_Mp9@4020_d N_OUT8_Mp9@4020_g N_VDD_Mp9@4020_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4019 N_OUT9_Mn9@4019_d N_OUT8_Mn9@4019_g N_VSS_Mn9@4019_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4018 N_OUT9_Mn9@4018_d N_OUT8_Mn9@4018_g N_VSS_Mn9@4018_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4019 N_OUT9_Mp9@4019_d N_OUT8_Mp9@4019_g N_VDD_Mp9@4019_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4018 N_OUT9_Mp9@4018_d N_OUT8_Mp9@4018_g N_VDD_Mp9@4018_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4017 N_OUT9_Mn9@4017_d N_OUT8_Mn9@4017_g N_VSS_Mn9@4017_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4016 N_OUT9_Mn9@4016_d N_OUT8_Mn9@4016_g N_VSS_Mn9@4016_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4017 N_OUT9_Mp9@4017_d N_OUT8_Mp9@4017_g N_VDD_Mp9@4017_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4016 N_OUT9_Mp9@4016_d N_OUT8_Mp9@4016_g N_VDD_Mp9@4016_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4015 N_OUT9_Mn9@4015_d N_OUT8_Mn9@4015_g N_VSS_Mn9@4015_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4014 N_OUT9_Mn9@4014_d N_OUT8_Mn9@4014_g N_VSS_Mn9@4014_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4015 N_OUT9_Mp9@4015_d N_OUT8_Mp9@4015_g N_VDD_Mp9@4015_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4014 N_OUT9_Mp9@4014_d N_OUT8_Mp9@4014_g N_VDD_Mp9@4014_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4013 N_OUT9_Mn9@4013_d N_OUT8_Mn9@4013_g N_VSS_Mn9@4013_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4012 N_OUT9_Mn9@4012_d N_OUT8_Mn9@4012_g N_VSS_Mn9@4012_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4013 N_OUT9_Mp9@4013_d N_OUT8_Mp9@4013_g N_VDD_Mp9@4013_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4012 N_OUT9_Mp9@4012_d N_OUT8_Mp9@4012_g N_VDD_Mp9@4012_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4011 N_OUT9_Mn9@4011_d N_OUT8_Mn9@4011_g N_VSS_Mn9@4011_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4010 N_OUT9_Mn9@4010_d N_OUT8_Mn9@4010_g N_VSS_Mn9@4010_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4011 N_OUT9_Mp9@4011_d N_OUT8_Mp9@4011_g N_VDD_Mp9@4011_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4010 N_OUT9_Mp9@4010_d N_OUT8_Mp9@4010_g N_VDD_Mp9@4010_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4009 N_OUT9_Mn9@4009_d N_OUT8_Mn9@4009_g N_VSS_Mn9@4009_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4008 N_OUT9_Mn9@4008_d N_OUT8_Mn9@4008_g N_VSS_Mn9@4008_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4009 N_OUT9_Mp9@4009_d N_OUT8_Mp9@4009_g N_VDD_Mp9@4009_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4008 N_OUT9_Mp9@4008_d N_OUT8_Mp9@4008_g N_VDD_Mp9@4008_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4007 N_OUT9_Mn9@4007_d N_OUT8_Mn9@4007_g N_VSS_Mn9@4007_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4006 N_OUT9_Mn9@4006_d N_OUT8_Mn9@4006_g N_VSS_Mn9@4006_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4007 N_OUT9_Mp9@4007_d N_OUT8_Mp9@4007_g N_VDD_Mp9@4007_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4006 N_OUT9_Mp9@4006_d N_OUT8_Mp9@4006_g N_VDD_Mp9@4006_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4005 N_OUT9_Mn9@4005_d N_OUT8_Mn9@4005_g N_VSS_Mn9@4005_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4004 N_OUT9_Mn9@4004_d N_OUT8_Mn9@4004_g N_VSS_Mn9@4004_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4005 N_OUT9_Mp9@4005_d N_OUT8_Mp9@4005_g N_VDD_Mp9@4005_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4004 N_OUT9_Mp9@4004_d N_OUT8_Mp9@4004_g N_VDD_Mp9@4004_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4003 N_OUT9_Mn9@4003_d N_OUT8_Mn9@4003_g N_VSS_Mn9@4003_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4002 N_OUT9_Mn9@4002_d N_OUT8_Mn9@4002_g N_VSS_Mn9@4002_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4003 N_OUT9_Mp9@4003_d N_OUT8_Mp9@4003_g N_VDD_Mp9@4003_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4002 N_OUT9_Mp9@4002_d N_OUT8_Mp9@4002_g N_VDD_Mp9@4002_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@4001 N_OUT9_Mn9@4001_d N_OUT8_Mn9@4001_g N_VSS_Mn9@4001_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4000 N_OUT9_Mn9@4000_d N_OUT8_Mn9@4000_g N_VSS_Mn9@4000_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@4001 N_OUT9_Mp9@4001_d N_OUT8_Mp9@4001_g N_VDD_Mp9@4001_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4000 N_OUT9_Mp9@4000_d N_OUT8_Mp9@4000_g N_VDD_Mp9@4000_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3999 N_OUT9_Mn9@3999_d N_OUT8_Mn9@3999_g N_VSS_Mn9@3999_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3998 N_OUT9_Mn9@3998_d N_OUT8_Mn9@3998_g N_VSS_Mn9@3998_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3999 N_OUT9_Mp9@3999_d N_OUT8_Mp9@3999_g N_VDD_Mp9@3999_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3998 N_OUT9_Mp9@3998_d N_OUT8_Mp9@3998_g N_VDD_Mp9@3998_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3997 N_OUT9_Mn9@3997_d N_OUT8_Mn9@3997_g N_VSS_Mn9@3997_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3996 N_OUT9_Mn9@3996_d N_OUT8_Mn9@3996_g N_VSS_Mn9@3996_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3997 N_OUT9_Mp9@3997_d N_OUT8_Mp9@3997_g N_VDD_Mp9@3997_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3996 N_OUT9_Mp9@3996_d N_OUT8_Mp9@3996_g N_VDD_Mp9@3996_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3995 N_OUT9_Mn9@3995_d N_OUT8_Mn9@3995_g N_VSS_Mn9@3995_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3994 N_OUT9_Mn9@3994_d N_OUT8_Mn9@3994_g N_VSS_Mn9@3994_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3995 N_OUT9_Mp9@3995_d N_OUT8_Mp9@3995_g N_VDD_Mp9@3995_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3994 N_OUT9_Mp9@3994_d N_OUT8_Mp9@3994_g N_VDD_Mp9@3994_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3993 N_OUT9_Mn9@3993_d N_OUT8_Mn9@3993_g N_VSS_Mn9@3993_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3992 N_OUT9_Mn9@3992_d N_OUT8_Mn9@3992_g N_VSS_Mn9@3992_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3993 N_OUT9_Mp9@3993_d N_OUT8_Mp9@3993_g N_VDD_Mp9@3993_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3992 N_OUT9_Mp9@3992_d N_OUT8_Mp9@3992_g N_VDD_Mp9@3992_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3991 N_OUT9_Mn9@3991_d N_OUT8_Mn9@3991_g N_VSS_Mn9@3991_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3990 N_OUT9_Mn9@3990_d N_OUT8_Mn9@3990_g N_VSS_Mn9@3990_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3991 N_OUT9_Mp9@3991_d N_OUT8_Mp9@3991_g N_VDD_Mp9@3991_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3990 N_OUT9_Mp9@3990_d N_OUT8_Mp9@3990_g N_VDD_Mp9@3990_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3989 N_OUT9_Mn9@3989_d N_OUT8_Mn9@3989_g N_VSS_Mn9@3989_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3988 N_OUT9_Mn9@3988_d N_OUT8_Mn9@3988_g N_VSS_Mn9@3988_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3989 N_OUT9_Mp9@3989_d N_OUT8_Mp9@3989_g N_VDD_Mp9@3989_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3988 N_OUT9_Mp9@3988_d N_OUT8_Mp9@3988_g N_VDD_Mp9@3988_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3987 N_OUT9_Mn9@3987_d N_OUT8_Mn9@3987_g N_VSS_Mn9@3987_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3986 N_OUT9_Mn9@3986_d N_OUT8_Mn9@3986_g N_VSS_Mn9@3986_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3987 N_OUT9_Mp9@3987_d N_OUT8_Mp9@3987_g N_VDD_Mp9@3987_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3986 N_OUT9_Mp9@3986_d N_OUT8_Mp9@3986_g N_VDD_Mp9@3986_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3985 N_OUT9_Mn9@3985_d N_OUT8_Mn9@3985_g N_VSS_Mn9@3985_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3984 N_OUT9_Mn9@3984_d N_OUT8_Mn9@3984_g N_VSS_Mn9@3984_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3985 N_OUT9_Mp9@3985_d N_OUT8_Mp9@3985_g N_VDD_Mp9@3985_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3984 N_OUT9_Mp9@3984_d N_OUT8_Mp9@3984_g N_VDD_Mp9@3984_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3983 N_OUT9_Mn9@3983_d N_OUT8_Mn9@3983_g N_VSS_Mn9@3983_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3982 N_OUT9_Mn9@3982_d N_OUT8_Mn9@3982_g N_VSS_Mn9@3982_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3983 N_OUT9_Mp9@3983_d N_OUT8_Mp9@3983_g N_VDD_Mp9@3983_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3982 N_OUT9_Mp9@3982_d N_OUT8_Mp9@3982_g N_VDD_Mp9@3982_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3981 N_OUT9_Mn9@3981_d N_OUT8_Mn9@3981_g N_VSS_Mn9@3981_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3980 N_OUT9_Mn9@3980_d N_OUT8_Mn9@3980_g N_VSS_Mn9@3980_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3981 N_OUT9_Mp9@3981_d N_OUT8_Mp9@3981_g N_VDD_Mp9@3981_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3980 N_OUT9_Mp9@3980_d N_OUT8_Mp9@3980_g N_VDD_Mp9@3980_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3979 N_OUT9_Mn9@3979_d N_OUT8_Mn9@3979_g N_VSS_Mn9@3979_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3978 N_OUT9_Mn9@3978_d N_OUT8_Mn9@3978_g N_VSS_Mn9@3978_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3979 N_OUT9_Mp9@3979_d N_OUT8_Mp9@3979_g N_VDD_Mp9@3979_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3978 N_OUT9_Mp9@3978_d N_OUT8_Mp9@3978_g N_VDD_Mp9@3978_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3977 N_OUT9_Mn9@3977_d N_OUT8_Mn9@3977_g N_VSS_Mn9@3977_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3976 N_OUT9_Mn9@3976_d N_OUT8_Mn9@3976_g N_VSS_Mn9@3976_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3977 N_OUT9_Mp9@3977_d N_OUT8_Mp9@3977_g N_VDD_Mp9@3977_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3976 N_OUT9_Mp9@3976_d N_OUT8_Mp9@3976_g N_VDD_Mp9@3976_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3975 N_OUT9_Mn9@3975_d N_OUT8_Mn9@3975_g N_VSS_Mn9@3975_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3974 N_OUT9_Mn9@3974_d N_OUT8_Mn9@3974_g N_VSS_Mn9@3974_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3975 N_OUT9_Mp9@3975_d N_OUT8_Mp9@3975_g N_VDD_Mp9@3975_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3974 N_OUT9_Mp9@3974_d N_OUT8_Mp9@3974_g N_VDD_Mp9@3974_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3973 N_OUT9_Mn9@3973_d N_OUT8_Mn9@3973_g N_VSS_Mn9@3973_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3972 N_OUT9_Mn9@3972_d N_OUT8_Mn9@3972_g N_VSS_Mn9@3972_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3973 N_OUT9_Mp9@3973_d N_OUT8_Mp9@3973_g N_VDD_Mp9@3973_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3972 N_OUT9_Mp9@3972_d N_OUT8_Mp9@3972_g N_VDD_Mp9@3972_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3971 N_OUT9_Mn9@3971_d N_OUT8_Mn9@3971_g N_VSS_Mn9@3971_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3970 N_OUT9_Mn9@3970_d N_OUT8_Mn9@3970_g N_VSS_Mn9@3970_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3971 N_OUT9_Mp9@3971_d N_OUT8_Mp9@3971_g N_VDD_Mp9@3971_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3970 N_OUT9_Mp9@3970_d N_OUT8_Mp9@3970_g N_VDD_Mp9@3970_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3969 N_OUT9_Mn9@3969_d N_OUT8_Mn9@3969_g N_VSS_Mn9@3969_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3968 N_OUT9_Mn9@3968_d N_OUT8_Mn9@3968_g N_VSS_Mn9@3968_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3969 N_OUT9_Mp9@3969_d N_OUT8_Mp9@3969_g N_VDD_Mp9@3969_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3968 N_OUT9_Mp9@3968_d N_OUT8_Mp9@3968_g N_VDD_Mp9@3968_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3967 N_OUT9_Mn9@3967_d N_OUT8_Mn9@3967_g N_VSS_Mn9@3967_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3966 N_OUT9_Mn9@3966_d N_OUT8_Mn9@3966_g N_VSS_Mn9@3966_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3967 N_OUT9_Mp9@3967_d N_OUT8_Mp9@3967_g N_VDD_Mp9@3967_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3966 N_OUT9_Mp9@3966_d N_OUT8_Mp9@3966_g N_VDD_Mp9@3966_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3965 N_OUT9_Mn9@3965_d N_OUT8_Mn9@3965_g N_VSS_Mn9@3965_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3964 N_OUT9_Mn9@3964_d N_OUT8_Mn9@3964_g N_VSS_Mn9@3964_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3965 N_OUT9_Mp9@3965_d N_OUT8_Mp9@3965_g N_VDD_Mp9@3965_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3964 N_OUT9_Mp9@3964_d N_OUT8_Mp9@3964_g N_VDD_Mp9@3964_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3963 N_OUT9_Mn9@3963_d N_OUT8_Mn9@3963_g N_VSS_Mn9@3963_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3962 N_OUT9_Mn9@3962_d N_OUT8_Mn9@3962_g N_VSS_Mn9@3962_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3963 N_OUT9_Mp9@3963_d N_OUT8_Mp9@3963_g N_VDD_Mp9@3963_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3962 N_OUT9_Mp9@3962_d N_OUT8_Mp9@3962_g N_VDD_Mp9@3962_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3961 N_OUT9_Mn9@3961_d N_OUT8_Mn9@3961_g N_VSS_Mn9@3961_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3960 N_OUT9_Mn9@3960_d N_OUT8_Mn9@3960_g N_VSS_Mn9@3960_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3961 N_OUT9_Mp9@3961_d N_OUT8_Mp9@3961_g N_VDD_Mp9@3961_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3960 N_OUT9_Mp9@3960_d N_OUT8_Mp9@3960_g N_VDD_Mp9@3960_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3959 N_OUT9_Mn9@3959_d N_OUT8_Mn9@3959_g N_VSS_Mn9@3959_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3958 N_OUT9_Mn9@3958_d N_OUT8_Mn9@3958_g N_VSS_Mn9@3958_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3959 N_OUT9_Mp9@3959_d N_OUT8_Mp9@3959_g N_VDD_Mp9@3959_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3958 N_OUT9_Mp9@3958_d N_OUT8_Mp9@3958_g N_VDD_Mp9@3958_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3957 N_OUT9_Mn9@3957_d N_OUT8_Mn9@3957_g N_VSS_Mn9@3957_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3956 N_OUT9_Mn9@3956_d N_OUT8_Mn9@3956_g N_VSS_Mn9@3956_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3957 N_OUT9_Mp9@3957_d N_OUT8_Mp9@3957_g N_VDD_Mp9@3957_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3956 N_OUT9_Mp9@3956_d N_OUT8_Mp9@3956_g N_VDD_Mp9@3956_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3955 N_OUT9_Mn9@3955_d N_OUT8_Mn9@3955_g N_VSS_Mn9@3955_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3954 N_OUT9_Mn9@3954_d N_OUT8_Mn9@3954_g N_VSS_Mn9@3954_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3955 N_OUT9_Mp9@3955_d N_OUT8_Mp9@3955_g N_VDD_Mp9@3955_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3954 N_OUT9_Mp9@3954_d N_OUT8_Mp9@3954_g N_VDD_Mp9@3954_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3953 N_OUT9_Mn9@3953_d N_OUT8_Mn9@3953_g N_VSS_Mn9@3953_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3952 N_OUT9_Mn9@3952_d N_OUT8_Mn9@3952_g N_VSS_Mn9@3952_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3953 N_OUT9_Mp9@3953_d N_OUT8_Mp9@3953_g N_VDD_Mp9@3953_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3952 N_OUT9_Mp9@3952_d N_OUT8_Mp9@3952_g N_VDD_Mp9@3952_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3951 N_OUT9_Mn9@3951_d N_OUT8_Mn9@3951_g N_VSS_Mn9@3951_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3950 N_OUT9_Mn9@3950_d N_OUT8_Mn9@3950_g N_VSS_Mn9@3950_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3951 N_OUT9_Mp9@3951_d N_OUT8_Mp9@3951_g N_VDD_Mp9@3951_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3950 N_OUT9_Mp9@3950_d N_OUT8_Mp9@3950_g N_VDD_Mp9@3950_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3949 N_OUT9_Mn9@3949_d N_OUT8_Mn9@3949_g N_VSS_Mn9@3949_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3948 N_OUT9_Mn9@3948_d N_OUT8_Mn9@3948_g N_VSS_Mn9@3948_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3949 N_OUT9_Mp9@3949_d N_OUT8_Mp9@3949_g N_VDD_Mp9@3949_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3948 N_OUT9_Mp9@3948_d N_OUT8_Mp9@3948_g N_VDD_Mp9@3948_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3947 N_OUT9_Mn9@3947_d N_OUT8_Mn9@3947_g N_VSS_Mn9@3947_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3946 N_OUT9_Mn9@3946_d N_OUT8_Mn9@3946_g N_VSS_Mn9@3946_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3947 N_OUT9_Mp9@3947_d N_OUT8_Mp9@3947_g N_VDD_Mp9@3947_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3946 N_OUT9_Mp9@3946_d N_OUT8_Mp9@3946_g N_VDD_Mp9@3946_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3945 N_OUT9_Mn9@3945_d N_OUT8_Mn9@3945_g N_VSS_Mn9@3945_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3944 N_OUT9_Mn9@3944_d N_OUT8_Mn9@3944_g N_VSS_Mn9@3944_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3945 N_OUT9_Mp9@3945_d N_OUT8_Mp9@3945_g N_VDD_Mp9@3945_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3944 N_OUT9_Mp9@3944_d N_OUT8_Mp9@3944_g N_VDD_Mp9@3944_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3943 N_OUT9_Mn9@3943_d N_OUT8_Mn9@3943_g N_VSS_Mn9@3943_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3942 N_OUT9_Mn9@3942_d N_OUT8_Mn9@3942_g N_VSS_Mn9@3942_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3943 N_OUT9_Mp9@3943_d N_OUT8_Mp9@3943_g N_VDD_Mp9@3943_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3942 N_OUT9_Mp9@3942_d N_OUT8_Mp9@3942_g N_VDD_Mp9@3942_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3941 N_OUT9_Mn9@3941_d N_OUT8_Mn9@3941_g N_VSS_Mn9@3941_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3940 N_OUT9_Mn9@3940_d N_OUT8_Mn9@3940_g N_VSS_Mn9@3940_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3941 N_OUT9_Mp9@3941_d N_OUT8_Mp9@3941_g N_VDD_Mp9@3941_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3940 N_OUT9_Mp9@3940_d N_OUT8_Mp9@3940_g N_VDD_Mp9@3940_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3939 N_OUT9_Mn9@3939_d N_OUT8_Mn9@3939_g N_VSS_Mn9@3939_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3938 N_OUT9_Mn9@3938_d N_OUT8_Mn9@3938_g N_VSS_Mn9@3938_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3939 N_OUT9_Mp9@3939_d N_OUT8_Mp9@3939_g N_VDD_Mp9@3939_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3938 N_OUT9_Mp9@3938_d N_OUT8_Mp9@3938_g N_VDD_Mp9@3938_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3937 N_OUT9_Mn9@3937_d N_OUT8_Mn9@3937_g N_VSS_Mn9@3937_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3936 N_OUT9_Mn9@3936_d N_OUT8_Mn9@3936_g N_VSS_Mn9@3936_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3937 N_OUT9_Mp9@3937_d N_OUT8_Mp9@3937_g N_VDD_Mp9@3937_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3936 N_OUT9_Mp9@3936_d N_OUT8_Mp9@3936_g N_VDD_Mp9@3936_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3935 N_OUT9_Mn9@3935_d N_OUT8_Mn9@3935_g N_VSS_Mn9@3935_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3934 N_OUT9_Mn9@3934_d N_OUT8_Mn9@3934_g N_VSS_Mn9@3934_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3935 N_OUT9_Mp9@3935_d N_OUT8_Mp9@3935_g N_VDD_Mp9@3935_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3934 N_OUT9_Mp9@3934_d N_OUT8_Mp9@3934_g N_VDD_Mp9@3934_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3933 N_OUT9_Mn9@3933_d N_OUT8_Mn9@3933_g N_VSS_Mn9@3933_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3932 N_OUT9_Mn9@3932_d N_OUT8_Mn9@3932_g N_VSS_Mn9@3932_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3933 N_OUT9_Mp9@3933_d N_OUT8_Mp9@3933_g N_VDD_Mp9@3933_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3932 N_OUT9_Mp9@3932_d N_OUT8_Mp9@3932_g N_VDD_Mp9@3932_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3931 N_OUT9_Mn9@3931_d N_OUT8_Mn9@3931_g N_VSS_Mn9@3931_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3930 N_OUT9_Mn9@3930_d N_OUT8_Mn9@3930_g N_VSS_Mn9@3930_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3931 N_OUT9_Mp9@3931_d N_OUT8_Mp9@3931_g N_VDD_Mp9@3931_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3930 N_OUT9_Mp9@3930_d N_OUT8_Mp9@3930_g N_VDD_Mp9@3930_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3929 N_OUT9_Mn9@3929_d N_OUT8_Mn9@3929_g N_VSS_Mn9@3929_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3928 N_OUT9_Mn9@3928_d N_OUT8_Mn9@3928_g N_VSS_Mn9@3928_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3929 N_OUT9_Mp9@3929_d N_OUT8_Mp9@3929_g N_VDD_Mp9@3929_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3928 N_OUT9_Mp9@3928_d N_OUT8_Mp9@3928_g N_VDD_Mp9@3928_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3927 N_OUT9_Mn9@3927_d N_OUT8_Mn9@3927_g N_VSS_Mn9@3927_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3926 N_OUT9_Mn9@3926_d N_OUT8_Mn9@3926_g N_VSS_Mn9@3926_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3927 N_OUT9_Mp9@3927_d N_OUT8_Mp9@3927_g N_VDD_Mp9@3927_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3926 N_OUT9_Mp9@3926_d N_OUT8_Mp9@3926_g N_VDD_Mp9@3926_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3925 N_OUT9_Mn9@3925_d N_OUT8_Mn9@3925_g N_VSS_Mn9@3925_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3924 N_OUT9_Mn9@3924_d N_OUT8_Mn9@3924_g N_VSS_Mn9@3924_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3925 N_OUT9_Mp9@3925_d N_OUT8_Mp9@3925_g N_VDD_Mp9@3925_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3924 N_OUT9_Mp9@3924_d N_OUT8_Mp9@3924_g N_VDD_Mp9@3924_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3923 N_OUT9_Mn9@3923_d N_OUT8_Mn9@3923_g N_VSS_Mn9@3923_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3922 N_OUT9_Mn9@3922_d N_OUT8_Mn9@3922_g N_VSS_Mn9@3922_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3923 N_OUT9_Mp9@3923_d N_OUT8_Mp9@3923_g N_VDD_Mp9@3923_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3922 N_OUT9_Mp9@3922_d N_OUT8_Mp9@3922_g N_VDD_Mp9@3922_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3921 N_OUT9_Mn9@3921_d N_OUT8_Mn9@3921_g N_VSS_Mn9@3921_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3920 N_OUT9_Mn9@3920_d N_OUT8_Mn9@3920_g N_VSS_Mn9@3920_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3921 N_OUT9_Mp9@3921_d N_OUT8_Mp9@3921_g N_VDD_Mp9@3921_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3920 N_OUT9_Mp9@3920_d N_OUT8_Mp9@3920_g N_VDD_Mp9@3920_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3919 N_OUT9_Mn9@3919_d N_OUT8_Mn9@3919_g N_VSS_Mn9@3919_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3918 N_OUT9_Mn9@3918_d N_OUT8_Mn9@3918_g N_VSS_Mn9@3918_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3919 N_OUT9_Mp9@3919_d N_OUT8_Mp9@3919_g N_VDD_Mp9@3919_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3918 N_OUT9_Mp9@3918_d N_OUT8_Mp9@3918_g N_VDD_Mp9@3918_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3917 N_OUT9_Mn9@3917_d N_OUT8_Mn9@3917_g N_VSS_Mn9@3917_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3916 N_OUT9_Mn9@3916_d N_OUT8_Mn9@3916_g N_VSS_Mn9@3916_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3917 N_OUT9_Mp9@3917_d N_OUT8_Mp9@3917_g N_VDD_Mp9@3917_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3916 N_OUT9_Mp9@3916_d N_OUT8_Mp9@3916_g N_VDD_Mp9@3916_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3915 N_OUT9_Mn9@3915_d N_OUT8_Mn9@3915_g N_VSS_Mn9@3915_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3914 N_OUT9_Mn9@3914_d N_OUT8_Mn9@3914_g N_VSS_Mn9@3914_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3915 N_OUT9_Mp9@3915_d N_OUT8_Mp9@3915_g N_VDD_Mp9@3915_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3914 N_OUT9_Mp9@3914_d N_OUT8_Mp9@3914_g N_VDD_Mp9@3914_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3913 N_OUT9_Mn9@3913_d N_OUT8_Mn9@3913_g N_VSS_Mn9@3913_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3912 N_OUT9_Mn9@3912_d N_OUT8_Mn9@3912_g N_VSS_Mn9@3912_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3913 N_OUT9_Mp9@3913_d N_OUT8_Mp9@3913_g N_VDD_Mp9@3913_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3912 N_OUT9_Mp9@3912_d N_OUT8_Mp9@3912_g N_VDD_Mp9@3912_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3911 N_OUT9_Mn9@3911_d N_OUT8_Mn9@3911_g N_VSS_Mn9@3911_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3910 N_OUT9_Mn9@3910_d N_OUT8_Mn9@3910_g N_VSS_Mn9@3910_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3911 N_OUT9_Mp9@3911_d N_OUT8_Mp9@3911_g N_VDD_Mp9@3911_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3910 N_OUT9_Mp9@3910_d N_OUT8_Mp9@3910_g N_VDD_Mp9@3910_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3909 N_OUT9_Mn9@3909_d N_OUT8_Mn9@3909_g N_VSS_Mn9@3909_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3908 N_OUT9_Mn9@3908_d N_OUT8_Mn9@3908_g N_VSS_Mn9@3908_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3909 N_OUT9_Mp9@3909_d N_OUT8_Mp9@3909_g N_VDD_Mp9@3909_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3908 N_OUT9_Mp9@3908_d N_OUT8_Mp9@3908_g N_VDD_Mp9@3908_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3907 N_OUT9_Mn9@3907_d N_OUT8_Mn9@3907_g N_VSS_Mn9@3907_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3906 N_OUT9_Mn9@3906_d N_OUT8_Mn9@3906_g N_VSS_Mn9@3906_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3907 N_OUT9_Mp9@3907_d N_OUT8_Mp9@3907_g N_VDD_Mp9@3907_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3906 N_OUT9_Mp9@3906_d N_OUT8_Mp9@3906_g N_VDD_Mp9@3906_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3905 N_OUT9_Mn9@3905_d N_OUT8_Mn9@3905_g N_VSS_Mn9@3905_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3904 N_OUT9_Mn9@3904_d N_OUT8_Mn9@3904_g N_VSS_Mn9@3904_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3905 N_OUT9_Mp9@3905_d N_OUT8_Mp9@3905_g N_VDD_Mp9@3905_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3904 N_OUT9_Mp9@3904_d N_OUT8_Mp9@3904_g N_VDD_Mp9@3904_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3903 N_OUT9_Mn9@3903_d N_OUT8_Mn9@3903_g N_VSS_Mn9@3903_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3902 N_OUT9_Mn9@3902_d N_OUT8_Mn9@3902_g N_VSS_Mn9@3902_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3903 N_OUT9_Mp9@3903_d N_OUT8_Mp9@3903_g N_VDD_Mp9@3903_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3902 N_OUT9_Mp9@3902_d N_OUT8_Mp9@3902_g N_VDD_Mp9@3902_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3901 N_OUT9_Mn9@3901_d N_OUT8_Mn9@3901_g N_VSS_Mn9@3901_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3900 N_OUT9_Mn9@3900_d N_OUT8_Mn9@3900_g N_VSS_Mn9@3900_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3901 N_OUT9_Mp9@3901_d N_OUT8_Mp9@3901_g N_VDD_Mp9@3901_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3900 N_OUT9_Mp9@3900_d N_OUT8_Mp9@3900_g N_VDD_Mp9@3900_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3899 N_OUT9_Mn9@3899_d N_OUT8_Mn9@3899_g N_VSS_Mn9@3899_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3898 N_OUT9_Mn9@3898_d N_OUT8_Mn9@3898_g N_VSS_Mn9@3898_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3899 N_OUT9_Mp9@3899_d N_OUT8_Mp9@3899_g N_VDD_Mp9@3899_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3898 N_OUT9_Mp9@3898_d N_OUT8_Mp9@3898_g N_VDD_Mp9@3898_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3897 N_OUT9_Mn9@3897_d N_OUT8_Mn9@3897_g N_VSS_Mn9@3897_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3896 N_OUT9_Mn9@3896_d N_OUT8_Mn9@3896_g N_VSS_Mn9@3896_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3897 N_OUT9_Mp9@3897_d N_OUT8_Mp9@3897_g N_VDD_Mp9@3897_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3896 N_OUT9_Mp9@3896_d N_OUT8_Mp9@3896_g N_VDD_Mp9@3896_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3895 N_OUT9_Mn9@3895_d N_OUT8_Mn9@3895_g N_VSS_Mn9@3895_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3894 N_OUT9_Mn9@3894_d N_OUT8_Mn9@3894_g N_VSS_Mn9@3894_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3895 N_OUT9_Mp9@3895_d N_OUT8_Mp9@3895_g N_VDD_Mp9@3895_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3894 N_OUT9_Mp9@3894_d N_OUT8_Mp9@3894_g N_VDD_Mp9@3894_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3893 N_OUT9_Mn9@3893_d N_OUT8_Mn9@3893_g N_VSS_Mn9@3893_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3892 N_OUT9_Mn9@3892_d N_OUT8_Mn9@3892_g N_VSS_Mn9@3892_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3893 N_OUT9_Mp9@3893_d N_OUT8_Mp9@3893_g N_VDD_Mp9@3893_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3892 N_OUT9_Mp9@3892_d N_OUT8_Mp9@3892_g N_VDD_Mp9@3892_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3891 N_OUT9_Mn9@3891_d N_OUT8_Mn9@3891_g N_VSS_Mn9@3891_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3890 N_OUT9_Mn9@3890_d N_OUT8_Mn9@3890_g N_VSS_Mn9@3890_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3891 N_OUT9_Mp9@3891_d N_OUT8_Mp9@3891_g N_VDD_Mp9@3891_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3890 N_OUT9_Mp9@3890_d N_OUT8_Mp9@3890_g N_VDD_Mp9@3890_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3889 N_OUT9_Mn9@3889_d N_OUT8_Mn9@3889_g N_VSS_Mn9@3889_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3888 N_OUT9_Mn9@3888_d N_OUT8_Mn9@3888_g N_VSS_Mn9@3888_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3889 N_OUT9_Mp9@3889_d N_OUT8_Mp9@3889_g N_VDD_Mp9@3889_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3888 N_OUT9_Mp9@3888_d N_OUT8_Mp9@3888_g N_VDD_Mp9@3888_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3887 N_OUT9_Mn9@3887_d N_OUT8_Mn9@3887_g N_VSS_Mn9@3887_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3886 N_OUT9_Mn9@3886_d N_OUT8_Mn9@3886_g N_VSS_Mn9@3886_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3887 N_OUT9_Mp9@3887_d N_OUT8_Mp9@3887_g N_VDD_Mp9@3887_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3886 N_OUT9_Mp9@3886_d N_OUT8_Mp9@3886_g N_VDD_Mp9@3886_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3885 N_OUT9_Mn9@3885_d N_OUT8_Mn9@3885_g N_VSS_Mn9@3885_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3884 N_OUT9_Mn9@3884_d N_OUT8_Mn9@3884_g N_VSS_Mn9@3884_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3885 N_OUT9_Mp9@3885_d N_OUT8_Mp9@3885_g N_VDD_Mp9@3885_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3884 N_OUT9_Mp9@3884_d N_OUT8_Mp9@3884_g N_VDD_Mp9@3884_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3883 N_OUT9_Mn9@3883_d N_OUT8_Mn9@3883_g N_VSS_Mn9@3883_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3882 N_OUT9_Mn9@3882_d N_OUT8_Mn9@3882_g N_VSS_Mn9@3882_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3883 N_OUT9_Mp9@3883_d N_OUT8_Mp9@3883_g N_VDD_Mp9@3883_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3882 N_OUT9_Mp9@3882_d N_OUT8_Mp9@3882_g N_VDD_Mp9@3882_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3881 N_OUT9_Mn9@3881_d N_OUT8_Mn9@3881_g N_VSS_Mn9@3881_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3880 N_OUT9_Mn9@3880_d N_OUT8_Mn9@3880_g N_VSS_Mn9@3880_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3881 N_OUT9_Mp9@3881_d N_OUT8_Mp9@3881_g N_VDD_Mp9@3881_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3880 N_OUT9_Mp9@3880_d N_OUT8_Mp9@3880_g N_VDD_Mp9@3880_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3879 N_OUT9_Mn9@3879_d N_OUT8_Mn9@3879_g N_VSS_Mn9@3879_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3878 N_OUT9_Mn9@3878_d N_OUT8_Mn9@3878_g N_VSS_Mn9@3878_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3879 N_OUT9_Mp9@3879_d N_OUT8_Mp9@3879_g N_VDD_Mp9@3879_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3878 N_OUT9_Mp9@3878_d N_OUT8_Mp9@3878_g N_VDD_Mp9@3878_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3877 N_OUT9_Mn9@3877_d N_OUT8_Mn9@3877_g N_VSS_Mn9@3877_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3876 N_OUT9_Mn9@3876_d N_OUT8_Mn9@3876_g N_VSS_Mn9@3876_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3877 N_OUT9_Mp9@3877_d N_OUT8_Mp9@3877_g N_VDD_Mp9@3877_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3876 N_OUT9_Mp9@3876_d N_OUT8_Mp9@3876_g N_VDD_Mp9@3876_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3875 N_OUT9_Mn9@3875_d N_OUT8_Mn9@3875_g N_VSS_Mn9@3875_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3874 N_OUT9_Mn9@3874_d N_OUT8_Mn9@3874_g N_VSS_Mn9@3874_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3875 N_OUT9_Mp9@3875_d N_OUT8_Mp9@3875_g N_VDD_Mp9@3875_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3874 N_OUT9_Mp9@3874_d N_OUT8_Mp9@3874_g N_VDD_Mp9@3874_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3873 N_OUT9_Mn9@3873_d N_OUT8_Mn9@3873_g N_VSS_Mn9@3873_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3872 N_OUT9_Mn9@3872_d N_OUT8_Mn9@3872_g N_VSS_Mn9@3872_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3873 N_OUT9_Mp9@3873_d N_OUT8_Mp9@3873_g N_VDD_Mp9@3873_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3872 N_OUT9_Mp9@3872_d N_OUT8_Mp9@3872_g N_VDD_Mp9@3872_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3871 N_OUT9_Mn9@3871_d N_OUT8_Mn9@3871_g N_VSS_Mn9@3871_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3870 N_OUT9_Mn9@3870_d N_OUT8_Mn9@3870_g N_VSS_Mn9@3870_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3871 N_OUT9_Mp9@3871_d N_OUT8_Mp9@3871_g N_VDD_Mp9@3871_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3870 N_OUT9_Mp9@3870_d N_OUT8_Mp9@3870_g N_VDD_Mp9@3870_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3869 N_OUT9_Mn9@3869_d N_OUT8_Mn9@3869_g N_VSS_Mn9@3869_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3868 N_OUT9_Mn9@3868_d N_OUT8_Mn9@3868_g N_VSS_Mn9@3868_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3869 N_OUT9_Mp9@3869_d N_OUT8_Mp9@3869_g N_VDD_Mp9@3869_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3868 N_OUT9_Mp9@3868_d N_OUT8_Mp9@3868_g N_VDD_Mp9@3868_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3867 N_OUT9_Mn9@3867_d N_OUT8_Mn9@3867_g N_VSS_Mn9@3867_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3866 N_OUT9_Mn9@3866_d N_OUT8_Mn9@3866_g N_VSS_Mn9@3866_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3867 N_OUT9_Mp9@3867_d N_OUT8_Mp9@3867_g N_VDD_Mp9@3867_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3866 N_OUT9_Mp9@3866_d N_OUT8_Mp9@3866_g N_VDD_Mp9@3866_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3865 N_OUT9_Mn9@3865_d N_OUT8_Mn9@3865_g N_VSS_Mn9@3865_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3864 N_OUT9_Mn9@3864_d N_OUT8_Mn9@3864_g N_VSS_Mn9@3864_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3865 N_OUT9_Mp9@3865_d N_OUT8_Mp9@3865_g N_VDD_Mp9@3865_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3864 N_OUT9_Mp9@3864_d N_OUT8_Mp9@3864_g N_VDD_Mp9@3864_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3863 N_OUT9_Mn9@3863_d N_OUT8_Mn9@3863_g N_VSS_Mn9@3863_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3862 N_OUT9_Mn9@3862_d N_OUT8_Mn9@3862_g N_VSS_Mn9@3862_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3863 N_OUT9_Mp9@3863_d N_OUT8_Mp9@3863_g N_VDD_Mp9@3863_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3862 N_OUT9_Mp9@3862_d N_OUT8_Mp9@3862_g N_VDD_Mp9@3862_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3861 N_OUT9_Mn9@3861_d N_OUT8_Mn9@3861_g N_VSS_Mn9@3861_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3860 N_OUT9_Mn9@3860_d N_OUT8_Mn9@3860_g N_VSS_Mn9@3860_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3861 N_OUT9_Mp9@3861_d N_OUT8_Mp9@3861_g N_VDD_Mp9@3861_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3860 N_OUT9_Mp9@3860_d N_OUT8_Mp9@3860_g N_VDD_Mp9@3860_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3859 N_OUT9_Mn9@3859_d N_OUT8_Mn9@3859_g N_VSS_Mn9@3859_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3858 N_OUT9_Mn9@3858_d N_OUT8_Mn9@3858_g N_VSS_Mn9@3858_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3859 N_OUT9_Mp9@3859_d N_OUT8_Mp9@3859_g N_VDD_Mp9@3859_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3858 N_OUT9_Mp9@3858_d N_OUT8_Mp9@3858_g N_VDD_Mp9@3858_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3857 N_OUT9_Mn9@3857_d N_OUT8_Mn9@3857_g N_VSS_Mn9@3857_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3856 N_OUT9_Mn9@3856_d N_OUT8_Mn9@3856_g N_VSS_Mn9@3856_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3857 N_OUT9_Mp9@3857_d N_OUT8_Mp9@3857_g N_VDD_Mp9@3857_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3856 N_OUT9_Mp9@3856_d N_OUT8_Mp9@3856_g N_VDD_Mp9@3856_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3855 N_OUT9_Mn9@3855_d N_OUT8_Mn9@3855_g N_VSS_Mn9@3855_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3854 N_OUT9_Mn9@3854_d N_OUT8_Mn9@3854_g N_VSS_Mn9@3854_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3855 N_OUT9_Mp9@3855_d N_OUT8_Mp9@3855_g N_VDD_Mp9@3855_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3854 N_OUT9_Mp9@3854_d N_OUT8_Mp9@3854_g N_VDD_Mp9@3854_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3853 N_OUT9_Mn9@3853_d N_OUT8_Mn9@3853_g N_VSS_Mn9@3853_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3852 N_OUT9_Mn9@3852_d N_OUT8_Mn9@3852_g N_VSS_Mn9@3852_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3853 N_OUT9_Mp9@3853_d N_OUT8_Mp9@3853_g N_VDD_Mp9@3853_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3852 N_OUT9_Mp9@3852_d N_OUT8_Mp9@3852_g N_VDD_Mp9@3852_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3851 N_OUT9_Mn9@3851_d N_OUT8_Mn9@3851_g N_VSS_Mn9@3851_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3850 N_OUT9_Mn9@3850_d N_OUT8_Mn9@3850_g N_VSS_Mn9@3850_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3851 N_OUT9_Mp9@3851_d N_OUT8_Mp9@3851_g N_VDD_Mp9@3851_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3850 N_OUT9_Mp9@3850_d N_OUT8_Mp9@3850_g N_VDD_Mp9@3850_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3849 N_OUT9_Mn9@3849_d N_OUT8_Mn9@3849_g N_VSS_Mn9@3849_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3848 N_OUT9_Mn9@3848_d N_OUT8_Mn9@3848_g N_VSS_Mn9@3848_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3849 N_OUT9_Mp9@3849_d N_OUT8_Mp9@3849_g N_VDD_Mp9@3849_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3848 N_OUT9_Mp9@3848_d N_OUT8_Mp9@3848_g N_VDD_Mp9@3848_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3847 N_OUT9_Mn9@3847_d N_OUT8_Mn9@3847_g N_VSS_Mn9@3847_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3846 N_OUT9_Mn9@3846_d N_OUT8_Mn9@3846_g N_VSS_Mn9@3846_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3847 N_OUT9_Mp9@3847_d N_OUT8_Mp9@3847_g N_VDD_Mp9@3847_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3846 N_OUT9_Mp9@3846_d N_OUT8_Mp9@3846_g N_VDD_Mp9@3846_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3845 N_OUT9_Mn9@3845_d N_OUT8_Mn9@3845_g N_VSS_Mn9@3845_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3844 N_OUT9_Mn9@3844_d N_OUT8_Mn9@3844_g N_VSS_Mn9@3844_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3845 N_OUT9_Mp9@3845_d N_OUT8_Mp9@3845_g N_VDD_Mp9@3845_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3844 N_OUT9_Mp9@3844_d N_OUT8_Mp9@3844_g N_VDD_Mp9@3844_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3843 N_OUT9_Mn9@3843_d N_OUT8_Mn9@3843_g N_VSS_Mn9@3843_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3842 N_OUT9_Mn9@3842_d N_OUT8_Mn9@3842_g N_VSS_Mn9@3842_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3843 N_OUT9_Mp9@3843_d N_OUT8_Mp9@3843_g N_VDD_Mp9@3843_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3842 N_OUT9_Mp9@3842_d N_OUT8_Mp9@3842_g N_VDD_Mp9@3842_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3841 N_OUT9_Mn9@3841_d N_OUT8_Mn9@3841_g N_VSS_Mn9@3841_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3840 N_OUT9_Mn9@3840_d N_OUT8_Mn9@3840_g N_VSS_Mn9@3840_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3841 N_OUT9_Mp9@3841_d N_OUT8_Mp9@3841_g N_VDD_Mp9@3841_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3840 N_OUT9_Mp9@3840_d N_OUT8_Mp9@3840_g N_VDD_Mp9@3840_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3839 N_OUT9_Mn9@3839_d N_OUT8_Mn9@3839_g N_VSS_Mn9@3839_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3838 N_OUT9_Mn9@3838_d N_OUT8_Mn9@3838_g N_VSS_Mn9@3838_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3839 N_OUT9_Mp9@3839_d N_OUT8_Mp9@3839_g N_VDD_Mp9@3839_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3838 N_OUT9_Mp9@3838_d N_OUT8_Mp9@3838_g N_VDD_Mp9@3838_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3837 N_OUT9_Mn9@3837_d N_OUT8_Mn9@3837_g N_VSS_Mn9@3837_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3836 N_OUT9_Mn9@3836_d N_OUT8_Mn9@3836_g N_VSS_Mn9@3836_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3837 N_OUT9_Mp9@3837_d N_OUT8_Mp9@3837_g N_VDD_Mp9@3837_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3836 N_OUT9_Mp9@3836_d N_OUT8_Mp9@3836_g N_VDD_Mp9@3836_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3835 N_OUT9_Mn9@3835_d N_OUT8_Mn9@3835_g N_VSS_Mn9@3835_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3834 N_OUT9_Mn9@3834_d N_OUT8_Mn9@3834_g N_VSS_Mn9@3834_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3835 N_OUT9_Mp9@3835_d N_OUT8_Mp9@3835_g N_VDD_Mp9@3835_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3834 N_OUT9_Mp9@3834_d N_OUT8_Mp9@3834_g N_VDD_Mp9@3834_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3833 N_OUT9_Mn9@3833_d N_OUT8_Mn9@3833_g N_VSS_Mn9@3833_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3832 N_OUT9_Mn9@3832_d N_OUT8_Mn9@3832_g N_VSS_Mn9@3832_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3833 N_OUT9_Mp9@3833_d N_OUT8_Mp9@3833_g N_VDD_Mp9@3833_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3832 N_OUT9_Mp9@3832_d N_OUT8_Mp9@3832_g N_VDD_Mp9@3832_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3831 N_OUT9_Mn9@3831_d N_OUT8_Mn9@3831_g N_VSS_Mn9@3831_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3830 N_OUT9_Mn9@3830_d N_OUT8_Mn9@3830_g N_VSS_Mn9@3830_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3831 N_OUT9_Mp9@3831_d N_OUT8_Mp9@3831_g N_VDD_Mp9@3831_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3830 N_OUT9_Mp9@3830_d N_OUT8_Mp9@3830_g N_VDD_Mp9@3830_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3829 N_OUT9_Mn9@3829_d N_OUT8_Mn9@3829_g N_VSS_Mn9@3829_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3828 N_OUT9_Mn9@3828_d N_OUT8_Mn9@3828_g N_VSS_Mn9@3828_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3829 N_OUT9_Mp9@3829_d N_OUT8_Mp9@3829_g N_VDD_Mp9@3829_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3828 N_OUT9_Mp9@3828_d N_OUT8_Mp9@3828_g N_VDD_Mp9@3828_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3827 N_OUT9_Mn9@3827_d N_OUT8_Mn9@3827_g N_VSS_Mn9@3827_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3826 N_OUT9_Mn9@3826_d N_OUT8_Mn9@3826_g N_VSS_Mn9@3826_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3827 N_OUT9_Mp9@3827_d N_OUT8_Mp9@3827_g N_VDD_Mp9@3827_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3826 N_OUT9_Mp9@3826_d N_OUT8_Mp9@3826_g N_VDD_Mp9@3826_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3825 N_OUT9_Mn9@3825_d N_OUT8_Mn9@3825_g N_VSS_Mn9@3825_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3824 N_OUT9_Mn9@3824_d N_OUT8_Mn9@3824_g N_VSS_Mn9@3824_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3825 N_OUT9_Mp9@3825_d N_OUT8_Mp9@3825_g N_VDD_Mp9@3825_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3824 N_OUT9_Mp9@3824_d N_OUT8_Mp9@3824_g N_VDD_Mp9@3824_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3823 N_OUT9_Mn9@3823_d N_OUT8_Mn9@3823_g N_VSS_Mn9@3823_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3822 N_OUT9_Mn9@3822_d N_OUT8_Mn9@3822_g N_VSS_Mn9@3822_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3823 N_OUT9_Mp9@3823_d N_OUT8_Mp9@3823_g N_VDD_Mp9@3823_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3822 N_OUT9_Mp9@3822_d N_OUT8_Mp9@3822_g N_VDD_Mp9@3822_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3821 N_OUT9_Mn9@3821_d N_OUT8_Mn9@3821_g N_VSS_Mn9@3821_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3820 N_OUT9_Mn9@3820_d N_OUT8_Mn9@3820_g N_VSS_Mn9@3820_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3821 N_OUT9_Mp9@3821_d N_OUT8_Mp9@3821_g N_VDD_Mp9@3821_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3820 N_OUT9_Mp9@3820_d N_OUT8_Mp9@3820_g N_VDD_Mp9@3820_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3819 N_OUT9_Mn9@3819_d N_OUT8_Mn9@3819_g N_VSS_Mn9@3819_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3818 N_OUT9_Mn9@3818_d N_OUT8_Mn9@3818_g N_VSS_Mn9@3818_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3819 N_OUT9_Mp9@3819_d N_OUT8_Mp9@3819_g N_VDD_Mp9@3819_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3818 N_OUT9_Mp9@3818_d N_OUT8_Mp9@3818_g N_VDD_Mp9@3818_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3817 N_OUT9_Mn9@3817_d N_OUT8_Mn9@3817_g N_VSS_Mn9@3817_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3816 N_OUT9_Mn9@3816_d N_OUT8_Mn9@3816_g N_VSS_Mn9@3816_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3817 N_OUT9_Mp9@3817_d N_OUT8_Mp9@3817_g N_VDD_Mp9@3817_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3816 N_OUT9_Mp9@3816_d N_OUT8_Mp9@3816_g N_VDD_Mp9@3816_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3815 N_OUT9_Mn9@3815_d N_OUT8_Mn9@3815_g N_VSS_Mn9@3815_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3814 N_OUT9_Mn9@3814_d N_OUT8_Mn9@3814_g N_VSS_Mn9@3814_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3815 N_OUT9_Mp9@3815_d N_OUT8_Mp9@3815_g N_VDD_Mp9@3815_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3814 N_OUT9_Mp9@3814_d N_OUT8_Mp9@3814_g N_VDD_Mp9@3814_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3813 N_OUT9_Mn9@3813_d N_OUT8_Mn9@3813_g N_VSS_Mn9@3813_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3812 N_OUT9_Mn9@3812_d N_OUT8_Mn9@3812_g N_VSS_Mn9@3812_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3813 N_OUT9_Mp9@3813_d N_OUT8_Mp9@3813_g N_VDD_Mp9@3813_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3812 N_OUT9_Mp9@3812_d N_OUT8_Mp9@3812_g N_VDD_Mp9@3812_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3811 N_OUT9_Mn9@3811_d N_OUT8_Mn9@3811_g N_VSS_Mn9@3811_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3810 N_OUT9_Mn9@3810_d N_OUT8_Mn9@3810_g N_VSS_Mn9@3810_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3811 N_OUT9_Mp9@3811_d N_OUT8_Mp9@3811_g N_VDD_Mp9@3811_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3810 N_OUT9_Mp9@3810_d N_OUT8_Mp9@3810_g N_VDD_Mp9@3810_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3809 N_OUT9_Mn9@3809_d N_OUT8_Mn9@3809_g N_VSS_Mn9@3809_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3808 N_OUT9_Mn9@3808_d N_OUT8_Mn9@3808_g N_VSS_Mn9@3808_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3809 N_OUT9_Mp9@3809_d N_OUT8_Mp9@3809_g N_VDD_Mp9@3809_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3808 N_OUT9_Mp9@3808_d N_OUT8_Mp9@3808_g N_VDD_Mp9@3808_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3807 N_OUT9_Mn9@3807_d N_OUT8_Mn9@3807_g N_VSS_Mn9@3807_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3806 N_OUT9_Mn9@3806_d N_OUT8_Mn9@3806_g N_VSS_Mn9@3806_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3807 N_OUT9_Mp9@3807_d N_OUT8_Mp9@3807_g N_VDD_Mp9@3807_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3806 N_OUT9_Mp9@3806_d N_OUT8_Mp9@3806_g N_VDD_Mp9@3806_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3805 N_OUT9_Mn9@3805_d N_OUT8_Mn9@3805_g N_VSS_Mn9@3805_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3804 N_OUT9_Mn9@3804_d N_OUT8_Mn9@3804_g N_VSS_Mn9@3804_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3805 N_OUT9_Mp9@3805_d N_OUT8_Mp9@3805_g N_VDD_Mp9@3805_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3804 N_OUT9_Mp9@3804_d N_OUT8_Mp9@3804_g N_VDD_Mp9@3804_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3803 N_OUT9_Mn9@3803_d N_OUT8_Mn9@3803_g N_VSS_Mn9@3803_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3802 N_OUT9_Mn9@3802_d N_OUT8_Mn9@3802_g N_VSS_Mn9@3802_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3803 N_OUT9_Mp9@3803_d N_OUT8_Mp9@3803_g N_VDD_Mp9@3803_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3802 N_OUT9_Mp9@3802_d N_OUT8_Mp9@3802_g N_VDD_Mp9@3802_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3801 N_OUT9_Mn9@3801_d N_OUT8_Mn9@3801_g N_VSS_Mn9@3801_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3800 N_OUT9_Mn9@3800_d N_OUT8_Mn9@3800_g N_VSS_Mn9@3800_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3801 N_OUT9_Mp9@3801_d N_OUT8_Mp9@3801_g N_VDD_Mp9@3801_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3800 N_OUT9_Mp9@3800_d N_OUT8_Mp9@3800_g N_VDD_Mp9@3800_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3799 N_OUT9_Mn9@3799_d N_OUT8_Mn9@3799_g N_VSS_Mn9@3799_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3798 N_OUT9_Mn9@3798_d N_OUT8_Mn9@3798_g N_VSS_Mn9@3798_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3799 N_OUT9_Mp9@3799_d N_OUT8_Mp9@3799_g N_VDD_Mp9@3799_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3798 N_OUT9_Mp9@3798_d N_OUT8_Mp9@3798_g N_VDD_Mp9@3798_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3797 N_OUT9_Mn9@3797_d N_OUT8_Mn9@3797_g N_VSS_Mn9@3797_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3796 N_OUT9_Mn9@3796_d N_OUT8_Mn9@3796_g N_VSS_Mn9@3796_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3797 N_OUT9_Mp9@3797_d N_OUT8_Mp9@3797_g N_VDD_Mp9@3797_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3796 N_OUT9_Mp9@3796_d N_OUT8_Mp9@3796_g N_VDD_Mp9@3796_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3795 N_OUT9_Mn9@3795_d N_OUT8_Mn9@3795_g N_VSS_Mn9@3795_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3794 N_OUT9_Mn9@3794_d N_OUT8_Mn9@3794_g N_VSS_Mn9@3794_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3795 N_OUT9_Mp9@3795_d N_OUT8_Mp9@3795_g N_VDD_Mp9@3795_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3794 N_OUT9_Mp9@3794_d N_OUT8_Mp9@3794_g N_VDD_Mp9@3794_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3793 N_OUT9_Mn9@3793_d N_OUT8_Mn9@3793_g N_VSS_Mn9@3793_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3792 N_OUT9_Mn9@3792_d N_OUT8_Mn9@3792_g N_VSS_Mn9@3792_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3793 N_OUT9_Mp9@3793_d N_OUT8_Mp9@3793_g N_VDD_Mp9@3793_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3792 N_OUT9_Mp9@3792_d N_OUT8_Mp9@3792_g N_VDD_Mp9@3792_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3791 N_OUT9_Mn9@3791_d N_OUT8_Mn9@3791_g N_VSS_Mn9@3791_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3790 N_OUT9_Mn9@3790_d N_OUT8_Mn9@3790_g N_VSS_Mn9@3790_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3791 N_OUT9_Mp9@3791_d N_OUT8_Mp9@3791_g N_VDD_Mp9@3791_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3790 N_OUT9_Mp9@3790_d N_OUT8_Mp9@3790_g N_VDD_Mp9@3790_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3789 N_OUT9_Mn9@3789_d N_OUT8_Mn9@3789_g N_VSS_Mn9@3789_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3788 N_OUT9_Mn9@3788_d N_OUT8_Mn9@3788_g N_VSS_Mn9@3788_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3789 N_OUT9_Mp9@3789_d N_OUT8_Mp9@3789_g N_VDD_Mp9@3789_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3788 N_OUT9_Mp9@3788_d N_OUT8_Mp9@3788_g N_VDD_Mp9@3788_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3787 N_OUT9_Mn9@3787_d N_OUT8_Mn9@3787_g N_VSS_Mn9@3787_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3786 N_OUT9_Mn9@3786_d N_OUT8_Mn9@3786_g N_VSS_Mn9@3786_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3787 N_OUT9_Mp9@3787_d N_OUT8_Mp9@3787_g N_VDD_Mp9@3787_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3786 N_OUT9_Mp9@3786_d N_OUT8_Mp9@3786_g N_VDD_Mp9@3786_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3785 N_OUT9_Mn9@3785_d N_OUT8_Mn9@3785_g N_VSS_Mn9@3785_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3784 N_OUT9_Mn9@3784_d N_OUT8_Mn9@3784_g N_VSS_Mn9@3784_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3785 N_OUT9_Mp9@3785_d N_OUT8_Mp9@3785_g N_VDD_Mp9@3785_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3784 N_OUT9_Mp9@3784_d N_OUT8_Mp9@3784_g N_VDD_Mp9@3784_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3783 N_OUT9_Mn9@3783_d N_OUT8_Mn9@3783_g N_VSS_Mn9@3783_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3782 N_OUT9_Mn9@3782_d N_OUT8_Mn9@3782_g N_VSS_Mn9@3782_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3783 N_OUT9_Mp9@3783_d N_OUT8_Mp9@3783_g N_VDD_Mp9@3783_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3782 N_OUT9_Mp9@3782_d N_OUT8_Mp9@3782_g N_VDD_Mp9@3782_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3781 N_OUT9_Mn9@3781_d N_OUT8_Mn9@3781_g N_VSS_Mn9@3781_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3780 N_OUT9_Mn9@3780_d N_OUT8_Mn9@3780_g N_VSS_Mn9@3780_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3781 N_OUT9_Mp9@3781_d N_OUT8_Mp9@3781_g N_VDD_Mp9@3781_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3780 N_OUT9_Mp9@3780_d N_OUT8_Mp9@3780_g N_VDD_Mp9@3780_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3779 N_OUT9_Mn9@3779_d N_OUT8_Mn9@3779_g N_VSS_Mn9@3779_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3778 N_OUT9_Mn9@3778_d N_OUT8_Mn9@3778_g N_VSS_Mn9@3778_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3779 N_OUT9_Mp9@3779_d N_OUT8_Mp9@3779_g N_VDD_Mp9@3779_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3778 N_OUT9_Mp9@3778_d N_OUT8_Mp9@3778_g N_VDD_Mp9@3778_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3777 N_OUT9_Mn9@3777_d N_OUT8_Mn9@3777_g N_VSS_Mn9@3777_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3776 N_OUT9_Mn9@3776_d N_OUT8_Mn9@3776_g N_VSS_Mn9@3776_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3777 N_OUT9_Mp9@3777_d N_OUT8_Mp9@3777_g N_VDD_Mp9@3777_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3776 N_OUT9_Mp9@3776_d N_OUT8_Mp9@3776_g N_VDD_Mp9@3776_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3775 N_OUT9_Mn9@3775_d N_OUT8_Mn9@3775_g N_VSS_Mn9@3775_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3774 N_OUT9_Mn9@3774_d N_OUT8_Mn9@3774_g N_VSS_Mn9@3774_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3775 N_OUT9_Mp9@3775_d N_OUT8_Mp9@3775_g N_VDD_Mp9@3775_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3774 N_OUT9_Mp9@3774_d N_OUT8_Mp9@3774_g N_VDD_Mp9@3774_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3773 N_OUT9_Mn9@3773_d N_OUT8_Mn9@3773_g N_VSS_Mn9@3773_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3772 N_OUT9_Mn9@3772_d N_OUT8_Mn9@3772_g N_VSS_Mn9@3772_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3773 N_OUT9_Mp9@3773_d N_OUT8_Mp9@3773_g N_VDD_Mp9@3773_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3772 N_OUT9_Mp9@3772_d N_OUT8_Mp9@3772_g N_VDD_Mp9@3772_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3771 N_OUT9_Mn9@3771_d N_OUT8_Mn9@3771_g N_VSS_Mn9@3771_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3770 N_OUT9_Mn9@3770_d N_OUT8_Mn9@3770_g N_VSS_Mn9@3770_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3771 N_OUT9_Mp9@3771_d N_OUT8_Mp9@3771_g N_VDD_Mp9@3771_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3770 N_OUT9_Mp9@3770_d N_OUT8_Mp9@3770_g N_VDD_Mp9@3770_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3769 N_OUT9_Mn9@3769_d N_OUT8_Mn9@3769_g N_VSS_Mn9@3769_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3768 N_OUT9_Mn9@3768_d N_OUT8_Mn9@3768_g N_VSS_Mn9@3768_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3769 N_OUT9_Mp9@3769_d N_OUT8_Mp9@3769_g N_VDD_Mp9@3769_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3768 N_OUT9_Mp9@3768_d N_OUT8_Mp9@3768_g N_VDD_Mp9@3768_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3767 N_OUT9_Mn9@3767_d N_OUT8_Mn9@3767_g N_VSS_Mn9@3767_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3766 N_OUT9_Mn9@3766_d N_OUT8_Mn9@3766_g N_VSS_Mn9@3766_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3767 N_OUT9_Mp9@3767_d N_OUT8_Mp9@3767_g N_VDD_Mp9@3767_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3766 N_OUT9_Mp9@3766_d N_OUT8_Mp9@3766_g N_VDD_Mp9@3766_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3765 N_OUT9_Mn9@3765_d N_OUT8_Mn9@3765_g N_VSS_Mn9@3765_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3764 N_OUT9_Mn9@3764_d N_OUT8_Mn9@3764_g N_VSS_Mn9@3764_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3765 N_OUT9_Mp9@3765_d N_OUT8_Mp9@3765_g N_VDD_Mp9@3765_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3764 N_OUT9_Mp9@3764_d N_OUT8_Mp9@3764_g N_VDD_Mp9@3764_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3763 N_OUT9_Mn9@3763_d N_OUT8_Mn9@3763_g N_VSS_Mn9@3763_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3762 N_OUT9_Mn9@3762_d N_OUT8_Mn9@3762_g N_VSS_Mn9@3762_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3763 N_OUT9_Mp9@3763_d N_OUT8_Mp9@3763_g N_VDD_Mp9@3763_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3762 N_OUT9_Mp9@3762_d N_OUT8_Mp9@3762_g N_VDD_Mp9@3762_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3761 N_OUT9_Mn9@3761_d N_OUT8_Mn9@3761_g N_VSS_Mn9@3761_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3760 N_OUT9_Mn9@3760_d N_OUT8_Mn9@3760_g N_VSS_Mn9@3760_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3761 N_OUT9_Mp9@3761_d N_OUT8_Mp9@3761_g N_VDD_Mp9@3761_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3760 N_OUT9_Mp9@3760_d N_OUT8_Mp9@3760_g N_VDD_Mp9@3760_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3759 N_OUT9_Mn9@3759_d N_OUT8_Mn9@3759_g N_VSS_Mn9@3759_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3758 N_OUT9_Mn9@3758_d N_OUT8_Mn9@3758_g N_VSS_Mn9@3758_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3759 N_OUT9_Mp9@3759_d N_OUT8_Mp9@3759_g N_VDD_Mp9@3759_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3758 N_OUT9_Mp9@3758_d N_OUT8_Mp9@3758_g N_VDD_Mp9@3758_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3757 N_OUT9_Mn9@3757_d N_OUT8_Mn9@3757_g N_VSS_Mn9@3757_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3756 N_OUT9_Mn9@3756_d N_OUT8_Mn9@3756_g N_VSS_Mn9@3756_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3757 N_OUT9_Mp9@3757_d N_OUT8_Mp9@3757_g N_VDD_Mp9@3757_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3756 N_OUT9_Mp9@3756_d N_OUT8_Mp9@3756_g N_VDD_Mp9@3756_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3755 N_OUT9_Mn9@3755_d N_OUT8_Mn9@3755_g N_VSS_Mn9@3755_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3754 N_OUT9_Mn9@3754_d N_OUT8_Mn9@3754_g N_VSS_Mn9@3754_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3755 N_OUT9_Mp9@3755_d N_OUT8_Mp9@3755_g N_VDD_Mp9@3755_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3754 N_OUT9_Mp9@3754_d N_OUT8_Mp9@3754_g N_VDD_Mp9@3754_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3753 N_OUT9_Mn9@3753_d N_OUT8_Mn9@3753_g N_VSS_Mn9@3753_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3752 N_OUT9_Mn9@3752_d N_OUT8_Mn9@3752_g N_VSS_Mn9@3752_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3753 N_OUT9_Mp9@3753_d N_OUT8_Mp9@3753_g N_VDD_Mp9@3753_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3752 N_OUT9_Mp9@3752_d N_OUT8_Mp9@3752_g N_VDD_Mp9@3752_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3751 N_OUT9_Mn9@3751_d N_OUT8_Mn9@3751_g N_VSS_Mn9@3751_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3750 N_OUT9_Mn9@3750_d N_OUT8_Mn9@3750_g N_VSS_Mn9@3750_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3751 N_OUT9_Mp9@3751_d N_OUT8_Mp9@3751_g N_VDD_Mp9@3751_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3750 N_OUT9_Mp9@3750_d N_OUT8_Mp9@3750_g N_VDD_Mp9@3750_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3749 N_OUT9_Mn9@3749_d N_OUT8_Mn9@3749_g N_VSS_Mn9@3749_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3748 N_OUT9_Mn9@3748_d N_OUT8_Mn9@3748_g N_VSS_Mn9@3748_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3749 N_OUT9_Mp9@3749_d N_OUT8_Mp9@3749_g N_VDD_Mp9@3749_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3748 N_OUT9_Mp9@3748_d N_OUT8_Mp9@3748_g N_VDD_Mp9@3748_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3747 N_OUT9_Mn9@3747_d N_OUT8_Mn9@3747_g N_VSS_Mn9@3747_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3746 N_OUT9_Mn9@3746_d N_OUT8_Mn9@3746_g N_VSS_Mn9@3746_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3747 N_OUT9_Mp9@3747_d N_OUT8_Mp9@3747_g N_VDD_Mp9@3747_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3746 N_OUT9_Mp9@3746_d N_OUT8_Mp9@3746_g N_VDD_Mp9@3746_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3745 N_OUT9_Mn9@3745_d N_OUT8_Mn9@3745_g N_VSS_Mn9@3745_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3744 N_OUT9_Mn9@3744_d N_OUT8_Mn9@3744_g N_VSS_Mn9@3744_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3745 N_OUT9_Mp9@3745_d N_OUT8_Mp9@3745_g N_VDD_Mp9@3745_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3744 N_OUT9_Mp9@3744_d N_OUT8_Mp9@3744_g N_VDD_Mp9@3744_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3743 N_OUT9_Mn9@3743_d N_OUT8_Mn9@3743_g N_VSS_Mn9@3743_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3742 N_OUT9_Mn9@3742_d N_OUT8_Mn9@3742_g N_VSS_Mn9@3742_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3743 N_OUT9_Mp9@3743_d N_OUT8_Mp9@3743_g N_VDD_Mp9@3743_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3742 N_OUT9_Mp9@3742_d N_OUT8_Mp9@3742_g N_VDD_Mp9@3742_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3741 N_OUT9_Mn9@3741_d N_OUT8_Mn9@3741_g N_VSS_Mn9@3741_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3740 N_OUT9_Mn9@3740_d N_OUT8_Mn9@3740_g N_VSS_Mn9@3740_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3741 N_OUT9_Mp9@3741_d N_OUT8_Mp9@3741_g N_VDD_Mp9@3741_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3740 N_OUT9_Mp9@3740_d N_OUT8_Mp9@3740_g N_VDD_Mp9@3740_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3739 N_OUT9_Mn9@3739_d N_OUT8_Mn9@3739_g N_VSS_Mn9@3739_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3738 N_OUT9_Mn9@3738_d N_OUT8_Mn9@3738_g N_VSS_Mn9@3738_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3739 N_OUT9_Mp9@3739_d N_OUT8_Mp9@3739_g N_VDD_Mp9@3739_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3738 N_OUT9_Mp9@3738_d N_OUT8_Mp9@3738_g N_VDD_Mp9@3738_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3737 N_OUT9_Mn9@3737_d N_OUT8_Mn9@3737_g N_VSS_Mn9@3737_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3736 N_OUT9_Mn9@3736_d N_OUT8_Mn9@3736_g N_VSS_Mn9@3736_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3737 N_OUT9_Mp9@3737_d N_OUT8_Mp9@3737_g N_VDD_Mp9@3737_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3736 N_OUT9_Mp9@3736_d N_OUT8_Mp9@3736_g N_VDD_Mp9@3736_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3735 N_OUT9_Mn9@3735_d N_OUT8_Mn9@3735_g N_VSS_Mn9@3735_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3734 N_OUT9_Mn9@3734_d N_OUT8_Mn9@3734_g N_VSS_Mn9@3734_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3735 N_OUT9_Mp9@3735_d N_OUT8_Mp9@3735_g N_VDD_Mp9@3735_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3734 N_OUT9_Mp9@3734_d N_OUT8_Mp9@3734_g N_VDD_Mp9@3734_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3733 N_OUT9_Mn9@3733_d N_OUT8_Mn9@3733_g N_VSS_Mn9@3733_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3732 N_OUT9_Mn9@3732_d N_OUT8_Mn9@3732_g N_VSS_Mn9@3732_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3733 N_OUT9_Mp9@3733_d N_OUT8_Mp9@3733_g N_VDD_Mp9@3733_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3732 N_OUT9_Mp9@3732_d N_OUT8_Mp9@3732_g N_VDD_Mp9@3732_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3731 N_OUT9_Mn9@3731_d N_OUT8_Mn9@3731_g N_VSS_Mn9@3731_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3730 N_OUT9_Mn9@3730_d N_OUT8_Mn9@3730_g N_VSS_Mn9@3730_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3731 N_OUT9_Mp9@3731_d N_OUT8_Mp9@3731_g N_VDD_Mp9@3731_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3730 N_OUT9_Mp9@3730_d N_OUT8_Mp9@3730_g N_VDD_Mp9@3730_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3729 N_OUT9_Mn9@3729_d N_OUT8_Mn9@3729_g N_VSS_Mn9@3729_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3728 N_OUT9_Mn9@3728_d N_OUT8_Mn9@3728_g N_VSS_Mn9@3728_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3729 N_OUT9_Mp9@3729_d N_OUT8_Mp9@3729_g N_VDD_Mp9@3729_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3728 N_OUT9_Mp9@3728_d N_OUT8_Mp9@3728_g N_VDD_Mp9@3728_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3727 N_OUT9_Mn9@3727_d N_OUT8_Mn9@3727_g N_VSS_Mn9@3727_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3726 N_OUT9_Mn9@3726_d N_OUT8_Mn9@3726_g N_VSS_Mn9@3726_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3727 N_OUT9_Mp9@3727_d N_OUT8_Mp9@3727_g N_VDD_Mp9@3727_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3726 N_OUT9_Mp9@3726_d N_OUT8_Mp9@3726_g N_VDD_Mp9@3726_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3725 N_OUT9_Mn9@3725_d N_OUT8_Mn9@3725_g N_VSS_Mn9@3725_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3724 N_OUT9_Mn9@3724_d N_OUT8_Mn9@3724_g N_VSS_Mn9@3724_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3725 N_OUT9_Mp9@3725_d N_OUT8_Mp9@3725_g N_VDD_Mp9@3725_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3724 N_OUT9_Mp9@3724_d N_OUT8_Mp9@3724_g N_VDD_Mp9@3724_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3723 N_OUT9_Mn9@3723_d N_OUT8_Mn9@3723_g N_VSS_Mn9@3723_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3722 N_OUT9_Mn9@3722_d N_OUT8_Mn9@3722_g N_VSS_Mn9@3722_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3723 N_OUT9_Mp9@3723_d N_OUT8_Mp9@3723_g N_VDD_Mp9@3723_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3722 N_OUT9_Mp9@3722_d N_OUT8_Mp9@3722_g N_VDD_Mp9@3722_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3721 N_OUT9_Mn9@3721_d N_OUT8_Mn9@3721_g N_VSS_Mn9@3721_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3720 N_OUT9_Mn9@3720_d N_OUT8_Mn9@3720_g N_VSS_Mn9@3720_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3721 N_OUT9_Mp9@3721_d N_OUT8_Mp9@3721_g N_VDD_Mp9@3721_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3720 N_OUT9_Mp9@3720_d N_OUT8_Mp9@3720_g N_VDD_Mp9@3720_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3719 N_OUT9_Mn9@3719_d N_OUT8_Mn9@3719_g N_VSS_Mn9@3719_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3718 N_OUT9_Mn9@3718_d N_OUT8_Mn9@3718_g N_VSS_Mn9@3718_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3719 N_OUT9_Mp9@3719_d N_OUT8_Mp9@3719_g N_VDD_Mp9@3719_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3718 N_OUT9_Mp9@3718_d N_OUT8_Mp9@3718_g N_VDD_Mp9@3718_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3717 N_OUT9_Mn9@3717_d N_OUT8_Mn9@3717_g N_VSS_Mn9@3717_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3716 N_OUT9_Mn9@3716_d N_OUT8_Mn9@3716_g N_VSS_Mn9@3716_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3717 N_OUT9_Mp9@3717_d N_OUT8_Mp9@3717_g N_VDD_Mp9@3717_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3716 N_OUT9_Mp9@3716_d N_OUT8_Mp9@3716_g N_VDD_Mp9@3716_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3715 N_OUT9_Mn9@3715_d N_OUT8_Mn9@3715_g N_VSS_Mn9@3715_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3714 N_OUT9_Mn9@3714_d N_OUT8_Mn9@3714_g N_VSS_Mn9@3714_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3715 N_OUT9_Mp9@3715_d N_OUT8_Mp9@3715_g N_VDD_Mp9@3715_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3714 N_OUT9_Mp9@3714_d N_OUT8_Mp9@3714_g N_VDD_Mp9@3714_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3713 N_OUT9_Mn9@3713_d N_OUT8_Mn9@3713_g N_VSS_Mn9@3713_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3712 N_OUT9_Mn9@3712_d N_OUT8_Mn9@3712_g N_VSS_Mn9@3712_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3713 N_OUT9_Mp9@3713_d N_OUT8_Mp9@3713_g N_VDD_Mp9@3713_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3712 N_OUT9_Mp9@3712_d N_OUT8_Mp9@3712_g N_VDD_Mp9@3712_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3711 N_OUT9_Mn9@3711_d N_OUT8_Mn9@3711_g N_VSS_Mn9@3711_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3710 N_OUT9_Mn9@3710_d N_OUT8_Mn9@3710_g N_VSS_Mn9@3710_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3711 N_OUT9_Mp9@3711_d N_OUT8_Mp9@3711_g N_VDD_Mp9@3711_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3710 N_OUT9_Mp9@3710_d N_OUT8_Mp9@3710_g N_VDD_Mp9@3710_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3709 N_OUT9_Mn9@3709_d N_OUT8_Mn9@3709_g N_VSS_Mn9@3709_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3708 N_OUT9_Mn9@3708_d N_OUT8_Mn9@3708_g N_VSS_Mn9@3708_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3709 N_OUT9_Mp9@3709_d N_OUT8_Mp9@3709_g N_VDD_Mp9@3709_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3708 N_OUT9_Mp9@3708_d N_OUT8_Mp9@3708_g N_VDD_Mp9@3708_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3707 N_OUT9_Mn9@3707_d N_OUT8_Mn9@3707_g N_VSS_Mn9@3707_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3706 N_OUT9_Mn9@3706_d N_OUT8_Mn9@3706_g N_VSS_Mn9@3706_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3707 N_OUT9_Mp9@3707_d N_OUT8_Mp9@3707_g N_VDD_Mp9@3707_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3706 N_OUT9_Mp9@3706_d N_OUT8_Mp9@3706_g N_VDD_Mp9@3706_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3705 N_OUT9_Mn9@3705_d N_OUT8_Mn9@3705_g N_VSS_Mn9@3705_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3704 N_OUT9_Mn9@3704_d N_OUT8_Mn9@3704_g N_VSS_Mn9@3704_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3705 N_OUT9_Mp9@3705_d N_OUT8_Mp9@3705_g N_VDD_Mp9@3705_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3704 N_OUT9_Mp9@3704_d N_OUT8_Mp9@3704_g N_VDD_Mp9@3704_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3703 N_OUT9_Mn9@3703_d N_OUT8_Mn9@3703_g N_VSS_Mn9@3703_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3702 N_OUT9_Mn9@3702_d N_OUT8_Mn9@3702_g N_VSS_Mn9@3702_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3703 N_OUT9_Mp9@3703_d N_OUT8_Mp9@3703_g N_VDD_Mp9@3703_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3702 N_OUT9_Mp9@3702_d N_OUT8_Mp9@3702_g N_VDD_Mp9@3702_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3701 N_OUT9_Mn9@3701_d N_OUT8_Mn9@3701_g N_VSS_Mn9@3701_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3700 N_OUT9_Mn9@3700_d N_OUT8_Mn9@3700_g N_VSS_Mn9@3700_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3701 N_OUT9_Mp9@3701_d N_OUT8_Mp9@3701_g N_VDD_Mp9@3701_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3700 N_OUT9_Mp9@3700_d N_OUT8_Mp9@3700_g N_VDD_Mp9@3700_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3699 N_OUT9_Mn9@3699_d N_OUT8_Mn9@3699_g N_VSS_Mn9@3699_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3698 N_OUT9_Mn9@3698_d N_OUT8_Mn9@3698_g N_VSS_Mn9@3698_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3699 N_OUT9_Mp9@3699_d N_OUT8_Mp9@3699_g N_VDD_Mp9@3699_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3698 N_OUT9_Mp9@3698_d N_OUT8_Mp9@3698_g N_VDD_Mp9@3698_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3697 N_OUT9_Mn9@3697_d N_OUT8_Mn9@3697_g N_VSS_Mn9@3697_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3696 N_OUT9_Mn9@3696_d N_OUT8_Mn9@3696_g N_VSS_Mn9@3696_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3697 N_OUT9_Mp9@3697_d N_OUT8_Mp9@3697_g N_VDD_Mp9@3697_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3696 N_OUT9_Mp9@3696_d N_OUT8_Mp9@3696_g N_VDD_Mp9@3696_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3695 N_OUT9_Mn9@3695_d N_OUT8_Mn9@3695_g N_VSS_Mn9@3695_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3694 N_OUT9_Mn9@3694_d N_OUT8_Mn9@3694_g N_VSS_Mn9@3694_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3695 N_OUT9_Mp9@3695_d N_OUT8_Mp9@3695_g N_VDD_Mp9@3695_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3694 N_OUT9_Mp9@3694_d N_OUT8_Mp9@3694_g N_VDD_Mp9@3694_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3693 N_OUT9_Mn9@3693_d N_OUT8_Mn9@3693_g N_VSS_Mn9@3693_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3692 N_OUT9_Mn9@3692_d N_OUT8_Mn9@3692_g N_VSS_Mn9@3692_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3693 N_OUT9_Mp9@3693_d N_OUT8_Mp9@3693_g N_VDD_Mp9@3693_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3692 N_OUT9_Mp9@3692_d N_OUT8_Mp9@3692_g N_VDD_Mp9@3692_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3691 N_OUT9_Mn9@3691_d N_OUT8_Mn9@3691_g N_VSS_Mn9@3691_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3690 N_OUT9_Mn9@3690_d N_OUT8_Mn9@3690_g N_VSS_Mn9@3690_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3691 N_OUT9_Mp9@3691_d N_OUT8_Mp9@3691_g N_VDD_Mp9@3691_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3690 N_OUT9_Mp9@3690_d N_OUT8_Mp9@3690_g N_VDD_Mp9@3690_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3689 N_OUT9_Mn9@3689_d N_OUT8_Mn9@3689_g N_VSS_Mn9@3689_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3688 N_OUT9_Mn9@3688_d N_OUT8_Mn9@3688_g N_VSS_Mn9@3688_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3689 N_OUT9_Mp9@3689_d N_OUT8_Mp9@3689_g N_VDD_Mp9@3689_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3688 N_OUT9_Mp9@3688_d N_OUT8_Mp9@3688_g N_VDD_Mp9@3688_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3687 N_OUT9_Mn9@3687_d N_OUT8_Mn9@3687_g N_VSS_Mn9@3687_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3686 N_OUT9_Mn9@3686_d N_OUT8_Mn9@3686_g N_VSS_Mn9@3686_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3687 N_OUT9_Mp9@3687_d N_OUT8_Mp9@3687_g N_VDD_Mp9@3687_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3686 N_OUT9_Mp9@3686_d N_OUT8_Mp9@3686_g N_VDD_Mp9@3686_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3685 N_OUT9_Mn9@3685_d N_OUT8_Mn9@3685_g N_VSS_Mn9@3685_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3684 N_OUT9_Mn9@3684_d N_OUT8_Mn9@3684_g N_VSS_Mn9@3684_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3685 N_OUT9_Mp9@3685_d N_OUT8_Mp9@3685_g N_VDD_Mp9@3685_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3684 N_OUT9_Mp9@3684_d N_OUT8_Mp9@3684_g N_VDD_Mp9@3684_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3683 N_OUT9_Mn9@3683_d N_OUT8_Mn9@3683_g N_VSS_Mn9@3683_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3682 N_OUT9_Mn9@3682_d N_OUT8_Mn9@3682_g N_VSS_Mn9@3682_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3683 N_OUT9_Mp9@3683_d N_OUT8_Mp9@3683_g N_VDD_Mp9@3683_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3682 N_OUT9_Mp9@3682_d N_OUT8_Mp9@3682_g N_VDD_Mp9@3682_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3681 N_OUT9_Mn9@3681_d N_OUT8_Mn9@3681_g N_VSS_Mn9@3681_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3680 N_OUT9_Mn9@3680_d N_OUT8_Mn9@3680_g N_VSS_Mn9@3680_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3681 N_OUT9_Mp9@3681_d N_OUT8_Mp9@3681_g N_VDD_Mp9@3681_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3680 N_OUT9_Mp9@3680_d N_OUT8_Mp9@3680_g N_VDD_Mp9@3680_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3679 N_OUT9_Mn9@3679_d N_OUT8_Mn9@3679_g N_VSS_Mn9@3679_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3678 N_OUT9_Mn9@3678_d N_OUT8_Mn9@3678_g N_VSS_Mn9@3678_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3679 N_OUT9_Mp9@3679_d N_OUT8_Mp9@3679_g N_VDD_Mp9@3679_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3678 N_OUT9_Mp9@3678_d N_OUT8_Mp9@3678_g N_VDD_Mp9@3678_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3677 N_OUT9_Mn9@3677_d N_OUT8_Mn9@3677_g N_VSS_Mn9@3677_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3676 N_OUT9_Mn9@3676_d N_OUT8_Mn9@3676_g N_VSS_Mn9@3676_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3677 N_OUT9_Mp9@3677_d N_OUT8_Mp9@3677_g N_VDD_Mp9@3677_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3676 N_OUT9_Mp9@3676_d N_OUT8_Mp9@3676_g N_VDD_Mp9@3676_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3675 N_OUT9_Mn9@3675_d N_OUT8_Mn9@3675_g N_VSS_Mn9@3675_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3674 N_OUT9_Mn9@3674_d N_OUT8_Mn9@3674_g N_VSS_Mn9@3674_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3675 N_OUT9_Mp9@3675_d N_OUT8_Mp9@3675_g N_VDD_Mp9@3675_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3674 N_OUT9_Mp9@3674_d N_OUT8_Mp9@3674_g N_VDD_Mp9@3674_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3673 N_OUT9_Mn9@3673_d N_OUT8_Mn9@3673_g N_VSS_Mn9@3673_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3672 N_OUT9_Mn9@3672_d N_OUT8_Mn9@3672_g N_VSS_Mn9@3672_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3673 N_OUT9_Mp9@3673_d N_OUT8_Mp9@3673_g N_VDD_Mp9@3673_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3672 N_OUT9_Mp9@3672_d N_OUT8_Mp9@3672_g N_VDD_Mp9@3672_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3671 N_OUT9_Mn9@3671_d N_OUT8_Mn9@3671_g N_VSS_Mn9@3671_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3670 N_OUT9_Mn9@3670_d N_OUT8_Mn9@3670_g N_VSS_Mn9@3670_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3671 N_OUT9_Mp9@3671_d N_OUT8_Mp9@3671_g N_VDD_Mp9@3671_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3670 N_OUT9_Mp9@3670_d N_OUT8_Mp9@3670_g N_VDD_Mp9@3670_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3669 N_OUT9_Mn9@3669_d N_OUT8_Mn9@3669_g N_VSS_Mn9@3669_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3668 N_OUT9_Mn9@3668_d N_OUT8_Mn9@3668_g N_VSS_Mn9@3668_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3669 N_OUT9_Mp9@3669_d N_OUT8_Mp9@3669_g N_VDD_Mp9@3669_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3668 N_OUT9_Mp9@3668_d N_OUT8_Mp9@3668_g N_VDD_Mp9@3668_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3667 N_OUT9_Mn9@3667_d N_OUT8_Mn9@3667_g N_VSS_Mn9@3667_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3666 N_OUT9_Mn9@3666_d N_OUT8_Mn9@3666_g N_VSS_Mn9@3666_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3667 N_OUT9_Mp9@3667_d N_OUT8_Mp9@3667_g N_VDD_Mp9@3667_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3666 N_OUT9_Mp9@3666_d N_OUT8_Mp9@3666_g N_VDD_Mp9@3666_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3665 N_OUT9_Mn9@3665_d N_OUT8_Mn9@3665_g N_VSS_Mn9@3665_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3664 N_OUT9_Mn9@3664_d N_OUT8_Mn9@3664_g N_VSS_Mn9@3664_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3665 N_OUT9_Mp9@3665_d N_OUT8_Mp9@3665_g N_VDD_Mp9@3665_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3664 N_OUT9_Mp9@3664_d N_OUT8_Mp9@3664_g N_VDD_Mp9@3664_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3663 N_OUT9_Mn9@3663_d N_OUT8_Mn9@3663_g N_VSS_Mn9@3663_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3662 N_OUT9_Mn9@3662_d N_OUT8_Mn9@3662_g N_VSS_Mn9@3662_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3663 N_OUT9_Mp9@3663_d N_OUT8_Mp9@3663_g N_VDD_Mp9@3663_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3662 N_OUT9_Mp9@3662_d N_OUT8_Mp9@3662_g N_VDD_Mp9@3662_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3661 N_OUT9_Mn9@3661_d N_OUT8_Mn9@3661_g N_VSS_Mn9@3661_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3660 N_OUT9_Mn9@3660_d N_OUT8_Mn9@3660_g N_VSS_Mn9@3660_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3661 N_OUT9_Mp9@3661_d N_OUT8_Mp9@3661_g N_VDD_Mp9@3661_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3660 N_OUT9_Mp9@3660_d N_OUT8_Mp9@3660_g N_VDD_Mp9@3660_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3659 N_OUT9_Mn9@3659_d N_OUT8_Mn9@3659_g N_VSS_Mn9@3659_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3658 N_OUT9_Mn9@3658_d N_OUT8_Mn9@3658_g N_VSS_Mn9@3658_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3659 N_OUT9_Mp9@3659_d N_OUT8_Mp9@3659_g N_VDD_Mp9@3659_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3658 N_OUT9_Mp9@3658_d N_OUT8_Mp9@3658_g N_VDD_Mp9@3658_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3657 N_OUT9_Mn9@3657_d N_OUT8_Mn9@3657_g N_VSS_Mn9@3657_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3656 N_OUT9_Mn9@3656_d N_OUT8_Mn9@3656_g N_VSS_Mn9@3656_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3657 N_OUT9_Mp9@3657_d N_OUT8_Mp9@3657_g N_VDD_Mp9@3657_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3656 N_OUT9_Mp9@3656_d N_OUT8_Mp9@3656_g N_VDD_Mp9@3656_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3655 N_OUT9_Mn9@3655_d N_OUT8_Mn9@3655_g N_VSS_Mn9@3655_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3654 N_OUT9_Mn9@3654_d N_OUT8_Mn9@3654_g N_VSS_Mn9@3654_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3655 N_OUT9_Mp9@3655_d N_OUT8_Mp9@3655_g N_VDD_Mp9@3655_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3654 N_OUT9_Mp9@3654_d N_OUT8_Mp9@3654_g N_VDD_Mp9@3654_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3653 N_OUT9_Mn9@3653_d N_OUT8_Mn9@3653_g N_VSS_Mn9@3653_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3652 N_OUT9_Mn9@3652_d N_OUT8_Mn9@3652_g N_VSS_Mn9@3652_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3653 N_OUT9_Mp9@3653_d N_OUT8_Mp9@3653_g N_VDD_Mp9@3653_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3652 N_OUT9_Mp9@3652_d N_OUT8_Mp9@3652_g N_VDD_Mp9@3652_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3651 N_OUT9_Mn9@3651_d N_OUT8_Mn9@3651_g N_VSS_Mn9@3651_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3650 N_OUT9_Mn9@3650_d N_OUT8_Mn9@3650_g N_VSS_Mn9@3650_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3651 N_OUT9_Mp9@3651_d N_OUT8_Mp9@3651_g N_VDD_Mp9@3651_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3650 N_OUT9_Mp9@3650_d N_OUT8_Mp9@3650_g N_VDD_Mp9@3650_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3649 N_OUT9_Mn9@3649_d N_OUT8_Mn9@3649_g N_VSS_Mn9@3649_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3648 N_OUT9_Mn9@3648_d N_OUT8_Mn9@3648_g N_VSS_Mn9@3648_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3649 N_OUT9_Mp9@3649_d N_OUT8_Mp9@3649_g N_VDD_Mp9@3649_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3648 N_OUT9_Mp9@3648_d N_OUT8_Mp9@3648_g N_VDD_Mp9@3648_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3647 N_OUT9_Mn9@3647_d N_OUT8_Mn9@3647_g N_VSS_Mn9@3647_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3646 N_OUT9_Mn9@3646_d N_OUT8_Mn9@3646_g N_VSS_Mn9@3646_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3647 N_OUT9_Mp9@3647_d N_OUT8_Mp9@3647_g N_VDD_Mp9@3647_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3646 N_OUT9_Mp9@3646_d N_OUT8_Mp9@3646_g N_VDD_Mp9@3646_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3645 N_OUT9_Mn9@3645_d N_OUT8_Mn9@3645_g N_VSS_Mn9@3645_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3644 N_OUT9_Mn9@3644_d N_OUT8_Mn9@3644_g N_VSS_Mn9@3644_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3645 N_OUT9_Mp9@3645_d N_OUT8_Mp9@3645_g N_VDD_Mp9@3645_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3644 N_OUT9_Mp9@3644_d N_OUT8_Mp9@3644_g N_VDD_Mp9@3644_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3643 N_OUT9_Mn9@3643_d N_OUT8_Mn9@3643_g N_VSS_Mn9@3643_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3642 N_OUT9_Mn9@3642_d N_OUT8_Mn9@3642_g N_VSS_Mn9@3642_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3643 N_OUT9_Mp9@3643_d N_OUT8_Mp9@3643_g N_VDD_Mp9@3643_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3642 N_OUT9_Mp9@3642_d N_OUT8_Mp9@3642_g N_VDD_Mp9@3642_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3641 N_OUT9_Mn9@3641_d N_OUT8_Mn9@3641_g N_VSS_Mn9@3641_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3640 N_OUT9_Mn9@3640_d N_OUT8_Mn9@3640_g N_VSS_Mn9@3640_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3641 N_OUT9_Mp9@3641_d N_OUT8_Mp9@3641_g N_VDD_Mp9@3641_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3640 N_OUT9_Mp9@3640_d N_OUT8_Mp9@3640_g N_VDD_Mp9@3640_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3639 N_OUT9_Mn9@3639_d N_OUT8_Mn9@3639_g N_VSS_Mn9@3639_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3638 N_OUT9_Mn9@3638_d N_OUT8_Mn9@3638_g N_VSS_Mn9@3638_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3639 N_OUT9_Mp9@3639_d N_OUT8_Mp9@3639_g N_VDD_Mp9@3639_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3638 N_OUT9_Mp9@3638_d N_OUT8_Mp9@3638_g N_VDD_Mp9@3638_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3637 N_OUT9_Mn9@3637_d N_OUT8_Mn9@3637_g N_VSS_Mn9@3637_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3636 N_OUT9_Mn9@3636_d N_OUT8_Mn9@3636_g N_VSS_Mn9@3636_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3637 N_OUT9_Mp9@3637_d N_OUT8_Mp9@3637_g N_VDD_Mp9@3637_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3636 N_OUT9_Mp9@3636_d N_OUT8_Mp9@3636_g N_VDD_Mp9@3636_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3635 N_OUT9_Mn9@3635_d N_OUT8_Mn9@3635_g N_VSS_Mn9@3635_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3634 N_OUT9_Mn9@3634_d N_OUT8_Mn9@3634_g N_VSS_Mn9@3634_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3635 N_OUT9_Mp9@3635_d N_OUT8_Mp9@3635_g N_VDD_Mp9@3635_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3634 N_OUT9_Mp9@3634_d N_OUT8_Mp9@3634_g N_VDD_Mp9@3634_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3633 N_OUT9_Mn9@3633_d N_OUT8_Mn9@3633_g N_VSS_Mn9@3633_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3632 N_OUT9_Mn9@3632_d N_OUT8_Mn9@3632_g N_VSS_Mn9@3632_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3633 N_OUT9_Mp9@3633_d N_OUT8_Mp9@3633_g N_VDD_Mp9@3633_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3632 N_OUT9_Mp9@3632_d N_OUT8_Mp9@3632_g N_VDD_Mp9@3632_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3631 N_OUT9_Mn9@3631_d N_OUT8_Mn9@3631_g N_VSS_Mn9@3631_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3630 N_OUT9_Mn9@3630_d N_OUT8_Mn9@3630_g N_VSS_Mn9@3630_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3631 N_OUT9_Mp9@3631_d N_OUT8_Mp9@3631_g N_VDD_Mp9@3631_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3630 N_OUT9_Mp9@3630_d N_OUT8_Mp9@3630_g N_VDD_Mp9@3630_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3629 N_OUT9_Mn9@3629_d N_OUT8_Mn9@3629_g N_VSS_Mn9@3629_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3628 N_OUT9_Mn9@3628_d N_OUT8_Mn9@3628_g N_VSS_Mn9@3628_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3629 N_OUT9_Mp9@3629_d N_OUT8_Mp9@3629_g N_VDD_Mp9@3629_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3628 N_OUT9_Mp9@3628_d N_OUT8_Mp9@3628_g N_VDD_Mp9@3628_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3627 N_OUT9_Mn9@3627_d N_OUT8_Mn9@3627_g N_VSS_Mn9@3627_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3626 N_OUT9_Mn9@3626_d N_OUT8_Mn9@3626_g N_VSS_Mn9@3626_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3627 N_OUT9_Mp9@3627_d N_OUT8_Mp9@3627_g N_VDD_Mp9@3627_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3626 N_OUT9_Mp9@3626_d N_OUT8_Mp9@3626_g N_VDD_Mp9@3626_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3625 N_OUT9_Mn9@3625_d N_OUT8_Mn9@3625_g N_VSS_Mn9@3625_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3624 N_OUT9_Mn9@3624_d N_OUT8_Mn9@3624_g N_VSS_Mn9@3624_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3625 N_OUT9_Mp9@3625_d N_OUT8_Mp9@3625_g N_VDD_Mp9@3625_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3624 N_OUT9_Mp9@3624_d N_OUT8_Mp9@3624_g N_VDD_Mp9@3624_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3623 N_OUT9_Mn9@3623_d N_OUT8_Mn9@3623_g N_VSS_Mn9@3623_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3622 N_OUT9_Mn9@3622_d N_OUT8_Mn9@3622_g N_VSS_Mn9@3622_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3623 N_OUT9_Mp9@3623_d N_OUT8_Mp9@3623_g N_VDD_Mp9@3623_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3622 N_OUT9_Mp9@3622_d N_OUT8_Mp9@3622_g N_VDD_Mp9@3622_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3621 N_OUT9_Mn9@3621_d N_OUT8_Mn9@3621_g N_VSS_Mn9@3621_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3620 N_OUT9_Mn9@3620_d N_OUT8_Mn9@3620_g N_VSS_Mn9@3620_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3621 N_OUT9_Mp9@3621_d N_OUT8_Mp9@3621_g N_VDD_Mp9@3621_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3620 N_OUT9_Mp9@3620_d N_OUT8_Mp9@3620_g N_VDD_Mp9@3620_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3619 N_OUT9_Mn9@3619_d N_OUT8_Mn9@3619_g N_VSS_Mn9@3619_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3618 N_OUT9_Mn9@3618_d N_OUT8_Mn9@3618_g N_VSS_Mn9@3618_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3619 N_OUT9_Mp9@3619_d N_OUT8_Mp9@3619_g N_VDD_Mp9@3619_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3618 N_OUT9_Mp9@3618_d N_OUT8_Mp9@3618_g N_VDD_Mp9@3618_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3617 N_OUT9_Mn9@3617_d N_OUT8_Mn9@3617_g N_VSS_Mn9@3617_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3616 N_OUT9_Mn9@3616_d N_OUT8_Mn9@3616_g N_VSS_Mn9@3616_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3617 N_OUT9_Mp9@3617_d N_OUT8_Mp9@3617_g N_VDD_Mp9@3617_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3616 N_OUT9_Mp9@3616_d N_OUT8_Mp9@3616_g N_VDD_Mp9@3616_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3615 N_OUT9_Mn9@3615_d N_OUT8_Mn9@3615_g N_VSS_Mn9@3615_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3614 N_OUT9_Mn9@3614_d N_OUT8_Mn9@3614_g N_VSS_Mn9@3614_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3615 N_OUT9_Mp9@3615_d N_OUT8_Mp9@3615_g N_VDD_Mp9@3615_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3614 N_OUT9_Mp9@3614_d N_OUT8_Mp9@3614_g N_VDD_Mp9@3614_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3613 N_OUT9_Mn9@3613_d N_OUT8_Mn9@3613_g N_VSS_Mn9@3613_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3612 N_OUT9_Mn9@3612_d N_OUT8_Mn9@3612_g N_VSS_Mn9@3612_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3613 N_OUT9_Mp9@3613_d N_OUT8_Mp9@3613_g N_VDD_Mp9@3613_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3612 N_OUT9_Mp9@3612_d N_OUT8_Mp9@3612_g N_VDD_Mp9@3612_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3611 N_OUT9_Mn9@3611_d N_OUT8_Mn9@3611_g N_VSS_Mn9@3611_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3610 N_OUT9_Mn9@3610_d N_OUT8_Mn9@3610_g N_VSS_Mn9@3610_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3611 N_OUT9_Mp9@3611_d N_OUT8_Mp9@3611_g N_VDD_Mp9@3611_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3610 N_OUT9_Mp9@3610_d N_OUT8_Mp9@3610_g N_VDD_Mp9@3610_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3609 N_OUT9_Mn9@3609_d N_OUT8_Mn9@3609_g N_VSS_Mn9@3609_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3608 N_OUT9_Mn9@3608_d N_OUT8_Mn9@3608_g N_VSS_Mn9@3608_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3609 N_OUT9_Mp9@3609_d N_OUT8_Mp9@3609_g N_VDD_Mp9@3609_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3608 N_OUT9_Mp9@3608_d N_OUT8_Mp9@3608_g N_VDD_Mp9@3608_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3607 N_OUT9_Mn9@3607_d N_OUT8_Mn9@3607_g N_VSS_Mn9@3607_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3606 N_OUT9_Mn9@3606_d N_OUT8_Mn9@3606_g N_VSS_Mn9@3606_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3607 N_OUT9_Mp9@3607_d N_OUT8_Mp9@3607_g N_VDD_Mp9@3607_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3606 N_OUT9_Mp9@3606_d N_OUT8_Mp9@3606_g N_VDD_Mp9@3606_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3605 N_OUT9_Mn9@3605_d N_OUT8_Mn9@3605_g N_VSS_Mn9@3605_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3604 N_OUT9_Mn9@3604_d N_OUT8_Mn9@3604_g N_VSS_Mn9@3604_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3605 N_OUT9_Mp9@3605_d N_OUT8_Mp9@3605_g N_VDD_Mp9@3605_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3604 N_OUT9_Mp9@3604_d N_OUT8_Mp9@3604_g N_VDD_Mp9@3604_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3603 N_OUT9_Mn9@3603_d N_OUT8_Mn9@3603_g N_VSS_Mn9@3603_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3602 N_OUT9_Mn9@3602_d N_OUT8_Mn9@3602_g N_VSS_Mn9@3602_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3603 N_OUT9_Mp9@3603_d N_OUT8_Mp9@3603_g N_VDD_Mp9@3603_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3602 N_OUT9_Mp9@3602_d N_OUT8_Mp9@3602_g N_VDD_Mp9@3602_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3601 N_OUT9_Mn9@3601_d N_OUT8_Mn9@3601_g N_VSS_Mn9@3601_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3600 N_OUT9_Mn9@3600_d N_OUT8_Mn9@3600_g N_VSS_Mn9@3600_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3601 N_OUT9_Mp9@3601_d N_OUT8_Mp9@3601_g N_VDD_Mp9@3601_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3600 N_OUT9_Mp9@3600_d N_OUT8_Mp9@3600_g N_VDD_Mp9@3600_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3599 N_OUT9_Mn9@3599_d N_OUT8_Mn9@3599_g N_VSS_Mn9@3599_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3598 N_OUT9_Mn9@3598_d N_OUT8_Mn9@3598_g N_VSS_Mn9@3598_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3599 N_OUT9_Mp9@3599_d N_OUT8_Mp9@3599_g N_VDD_Mp9@3599_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3598 N_OUT9_Mp9@3598_d N_OUT8_Mp9@3598_g N_VDD_Mp9@3598_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3597 N_OUT9_Mn9@3597_d N_OUT8_Mn9@3597_g N_VSS_Mn9@3597_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3596 N_OUT9_Mn9@3596_d N_OUT8_Mn9@3596_g N_VSS_Mn9@3596_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3597 N_OUT9_Mp9@3597_d N_OUT8_Mp9@3597_g N_VDD_Mp9@3597_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3596 N_OUT9_Mp9@3596_d N_OUT8_Mp9@3596_g N_VDD_Mp9@3596_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3595 N_OUT9_Mn9@3595_d N_OUT8_Mn9@3595_g N_VSS_Mn9@3595_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3594 N_OUT9_Mn9@3594_d N_OUT8_Mn9@3594_g N_VSS_Mn9@3594_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3595 N_OUT9_Mp9@3595_d N_OUT8_Mp9@3595_g N_VDD_Mp9@3595_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3594 N_OUT9_Mp9@3594_d N_OUT8_Mp9@3594_g N_VDD_Mp9@3594_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3593 N_OUT9_Mn9@3593_d N_OUT8_Mn9@3593_g N_VSS_Mn9@3593_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3592 N_OUT9_Mn9@3592_d N_OUT8_Mn9@3592_g N_VSS_Mn9@3592_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3593 N_OUT9_Mp9@3593_d N_OUT8_Mp9@3593_g N_VDD_Mp9@3593_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3592 N_OUT9_Mp9@3592_d N_OUT8_Mp9@3592_g N_VDD_Mp9@3592_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3591 N_OUT9_Mn9@3591_d N_OUT8_Mn9@3591_g N_VSS_Mn9@3591_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3590 N_OUT9_Mn9@3590_d N_OUT8_Mn9@3590_g N_VSS_Mn9@3590_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3591 N_OUT9_Mp9@3591_d N_OUT8_Mp9@3591_g N_VDD_Mp9@3591_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3590 N_OUT9_Mp9@3590_d N_OUT8_Mp9@3590_g N_VDD_Mp9@3590_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3589 N_OUT9_Mn9@3589_d N_OUT8_Mn9@3589_g N_VSS_Mn9@3589_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3588 N_OUT9_Mn9@3588_d N_OUT8_Mn9@3588_g N_VSS_Mn9@3588_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3589 N_OUT9_Mp9@3589_d N_OUT8_Mp9@3589_g N_VDD_Mp9@3589_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3588 N_OUT9_Mp9@3588_d N_OUT8_Mp9@3588_g N_VDD_Mp9@3588_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3587 N_OUT9_Mn9@3587_d N_OUT8_Mn9@3587_g N_VSS_Mn9@3587_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3586 N_OUT9_Mn9@3586_d N_OUT8_Mn9@3586_g N_VSS_Mn9@3586_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3587 N_OUT9_Mp9@3587_d N_OUT8_Mp9@3587_g N_VDD_Mp9@3587_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3586 N_OUT9_Mp9@3586_d N_OUT8_Mp9@3586_g N_VDD_Mp9@3586_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3585 N_OUT9_Mn9@3585_d N_OUT8_Mn9@3585_g N_VSS_Mn9@3585_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3584 N_OUT9_Mn9@3584_d N_OUT8_Mn9@3584_g N_VSS_Mn9@3584_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3585 N_OUT9_Mp9@3585_d N_OUT8_Mp9@3585_g N_VDD_Mp9@3585_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3584 N_OUT9_Mp9@3584_d N_OUT8_Mp9@3584_g N_VDD_Mp9@3584_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3583 N_OUT9_Mn9@3583_d N_OUT8_Mn9@3583_g N_VSS_Mn9@3583_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3582 N_OUT9_Mn9@3582_d N_OUT8_Mn9@3582_g N_VSS_Mn9@3582_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3583 N_OUT9_Mp9@3583_d N_OUT8_Mp9@3583_g N_VDD_Mp9@3583_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3582 N_OUT9_Mp9@3582_d N_OUT8_Mp9@3582_g N_VDD_Mp9@3582_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3581 N_OUT9_Mn9@3581_d N_OUT8_Mn9@3581_g N_VSS_Mn9@3581_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3580 N_OUT9_Mn9@3580_d N_OUT8_Mn9@3580_g N_VSS_Mn9@3580_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3581 N_OUT9_Mp9@3581_d N_OUT8_Mp9@3581_g N_VDD_Mp9@3581_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3580 N_OUT9_Mp9@3580_d N_OUT8_Mp9@3580_g N_VDD_Mp9@3580_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3579 N_OUT9_Mn9@3579_d N_OUT8_Mn9@3579_g N_VSS_Mn9@3579_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3578 N_OUT9_Mn9@3578_d N_OUT8_Mn9@3578_g N_VSS_Mn9@3578_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3579 N_OUT9_Mp9@3579_d N_OUT8_Mp9@3579_g N_VDD_Mp9@3579_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3578 N_OUT9_Mp9@3578_d N_OUT8_Mp9@3578_g N_VDD_Mp9@3578_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3577 N_OUT9_Mn9@3577_d N_OUT8_Mn9@3577_g N_VSS_Mn9@3577_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3576 N_OUT9_Mn9@3576_d N_OUT8_Mn9@3576_g N_VSS_Mn9@3576_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3577 N_OUT9_Mp9@3577_d N_OUT8_Mp9@3577_g N_VDD_Mp9@3577_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3576 N_OUT9_Mp9@3576_d N_OUT8_Mp9@3576_g N_VDD_Mp9@3576_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3575 N_OUT9_Mn9@3575_d N_OUT8_Mn9@3575_g N_VSS_Mn9@3575_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3574 N_OUT9_Mn9@3574_d N_OUT8_Mn9@3574_g N_VSS_Mn9@3574_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3575 N_OUT9_Mp9@3575_d N_OUT8_Mp9@3575_g N_VDD_Mp9@3575_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3574 N_OUT9_Mp9@3574_d N_OUT8_Mp9@3574_g N_VDD_Mp9@3574_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3573 N_OUT9_Mn9@3573_d N_OUT8_Mn9@3573_g N_VSS_Mn9@3573_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3572 N_OUT9_Mn9@3572_d N_OUT8_Mn9@3572_g N_VSS_Mn9@3572_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3573 N_OUT9_Mp9@3573_d N_OUT8_Mp9@3573_g N_VDD_Mp9@3573_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3572 N_OUT9_Mp9@3572_d N_OUT8_Mp9@3572_g N_VDD_Mp9@3572_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3571 N_OUT9_Mn9@3571_d N_OUT8_Mn9@3571_g N_VSS_Mn9@3571_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3570 N_OUT9_Mn9@3570_d N_OUT8_Mn9@3570_g N_VSS_Mn9@3570_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3571 N_OUT9_Mp9@3571_d N_OUT8_Mp9@3571_g N_VDD_Mp9@3571_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3570 N_OUT9_Mp9@3570_d N_OUT8_Mp9@3570_g N_VDD_Mp9@3570_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3569 N_OUT9_Mn9@3569_d N_OUT8_Mn9@3569_g N_VSS_Mn9@3569_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3568 N_OUT9_Mn9@3568_d N_OUT8_Mn9@3568_g N_VSS_Mn9@3568_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3569 N_OUT9_Mp9@3569_d N_OUT8_Mp9@3569_g N_VDD_Mp9@3569_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3568 N_OUT9_Mp9@3568_d N_OUT8_Mp9@3568_g N_VDD_Mp9@3568_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3567 N_OUT9_Mn9@3567_d N_OUT8_Mn9@3567_g N_VSS_Mn9@3567_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3566 N_OUT9_Mn9@3566_d N_OUT8_Mn9@3566_g N_VSS_Mn9@3566_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3567 N_OUT9_Mp9@3567_d N_OUT8_Mp9@3567_g N_VDD_Mp9@3567_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3566 N_OUT9_Mp9@3566_d N_OUT8_Mp9@3566_g N_VDD_Mp9@3566_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3565 N_OUT9_Mn9@3565_d N_OUT8_Mn9@3565_g N_VSS_Mn9@3565_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3564 N_OUT9_Mn9@3564_d N_OUT8_Mn9@3564_g N_VSS_Mn9@3564_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3565 N_OUT9_Mp9@3565_d N_OUT8_Mp9@3565_g N_VDD_Mp9@3565_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3564 N_OUT9_Mp9@3564_d N_OUT8_Mp9@3564_g N_VDD_Mp9@3564_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3563 N_OUT9_Mn9@3563_d N_OUT8_Mn9@3563_g N_VSS_Mn9@3563_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3562 N_OUT9_Mn9@3562_d N_OUT8_Mn9@3562_g N_VSS_Mn9@3562_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3563 N_OUT9_Mp9@3563_d N_OUT8_Mp9@3563_g N_VDD_Mp9@3563_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3562 N_OUT9_Mp9@3562_d N_OUT8_Mp9@3562_g N_VDD_Mp9@3562_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3561 N_OUT9_Mn9@3561_d N_OUT8_Mn9@3561_g N_VSS_Mn9@3561_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3560 N_OUT9_Mn9@3560_d N_OUT8_Mn9@3560_g N_VSS_Mn9@3560_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3561 N_OUT9_Mp9@3561_d N_OUT8_Mp9@3561_g N_VDD_Mp9@3561_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3560 N_OUT9_Mp9@3560_d N_OUT8_Mp9@3560_g N_VDD_Mp9@3560_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3559 N_OUT9_Mn9@3559_d N_OUT8_Mn9@3559_g N_VSS_Mn9@3559_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3558 N_OUT9_Mn9@3558_d N_OUT8_Mn9@3558_g N_VSS_Mn9@3558_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3559 N_OUT9_Mp9@3559_d N_OUT8_Mp9@3559_g N_VDD_Mp9@3559_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3558 N_OUT9_Mp9@3558_d N_OUT8_Mp9@3558_g N_VDD_Mp9@3558_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3557 N_OUT9_Mn9@3557_d N_OUT8_Mn9@3557_g N_VSS_Mn9@3557_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3556 N_OUT9_Mn9@3556_d N_OUT8_Mn9@3556_g N_VSS_Mn9@3556_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3557 N_OUT9_Mp9@3557_d N_OUT8_Mp9@3557_g N_VDD_Mp9@3557_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3556 N_OUT9_Mp9@3556_d N_OUT8_Mp9@3556_g N_VDD_Mp9@3556_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3555 N_OUT9_Mn9@3555_d N_OUT8_Mn9@3555_g N_VSS_Mn9@3555_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3554 N_OUT9_Mn9@3554_d N_OUT8_Mn9@3554_g N_VSS_Mn9@3554_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3555 N_OUT9_Mp9@3555_d N_OUT8_Mp9@3555_g N_VDD_Mp9@3555_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3554 N_OUT9_Mp9@3554_d N_OUT8_Mp9@3554_g N_VDD_Mp9@3554_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3553 N_OUT9_Mn9@3553_d N_OUT8_Mn9@3553_g N_VSS_Mn9@3553_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3552 N_OUT9_Mn9@3552_d N_OUT8_Mn9@3552_g N_VSS_Mn9@3552_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3553 N_OUT9_Mp9@3553_d N_OUT8_Mp9@3553_g N_VDD_Mp9@3553_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3552 N_OUT9_Mp9@3552_d N_OUT8_Mp9@3552_g N_VDD_Mp9@3552_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3551 N_OUT9_Mn9@3551_d N_OUT8_Mn9@3551_g N_VSS_Mn9@3551_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3550 N_OUT9_Mn9@3550_d N_OUT8_Mn9@3550_g N_VSS_Mn9@3550_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3551 N_OUT9_Mp9@3551_d N_OUT8_Mp9@3551_g N_VDD_Mp9@3551_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3550 N_OUT9_Mp9@3550_d N_OUT8_Mp9@3550_g N_VDD_Mp9@3550_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3549 N_OUT9_Mn9@3549_d N_OUT8_Mn9@3549_g N_VSS_Mn9@3549_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3548 N_OUT9_Mn9@3548_d N_OUT8_Mn9@3548_g N_VSS_Mn9@3548_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3549 N_OUT9_Mp9@3549_d N_OUT8_Mp9@3549_g N_VDD_Mp9@3549_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3548 N_OUT9_Mp9@3548_d N_OUT8_Mp9@3548_g N_VDD_Mp9@3548_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3547 N_OUT9_Mn9@3547_d N_OUT8_Mn9@3547_g N_VSS_Mn9@3547_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3546 N_OUT9_Mn9@3546_d N_OUT8_Mn9@3546_g N_VSS_Mn9@3546_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3547 N_OUT9_Mp9@3547_d N_OUT8_Mp9@3547_g N_VDD_Mp9@3547_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3546 N_OUT9_Mp9@3546_d N_OUT8_Mp9@3546_g N_VDD_Mp9@3546_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3545 N_OUT9_Mn9@3545_d N_OUT8_Mn9@3545_g N_VSS_Mn9@3545_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3544 N_OUT9_Mn9@3544_d N_OUT8_Mn9@3544_g N_VSS_Mn9@3544_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3545 N_OUT9_Mp9@3545_d N_OUT8_Mp9@3545_g N_VDD_Mp9@3545_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3544 N_OUT9_Mp9@3544_d N_OUT8_Mp9@3544_g N_VDD_Mp9@3544_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3543 N_OUT9_Mn9@3543_d N_OUT8_Mn9@3543_g N_VSS_Mn9@3543_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3542 N_OUT9_Mn9@3542_d N_OUT8_Mn9@3542_g N_VSS_Mn9@3542_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3543 N_OUT9_Mp9@3543_d N_OUT8_Mp9@3543_g N_VDD_Mp9@3543_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3542 N_OUT9_Mp9@3542_d N_OUT8_Mp9@3542_g N_VDD_Mp9@3542_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3541 N_OUT9_Mn9@3541_d N_OUT8_Mn9@3541_g N_VSS_Mn9@3541_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3540 N_OUT9_Mn9@3540_d N_OUT8_Mn9@3540_g N_VSS_Mn9@3540_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3541 N_OUT9_Mp9@3541_d N_OUT8_Mp9@3541_g N_VDD_Mp9@3541_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3540 N_OUT9_Mp9@3540_d N_OUT8_Mp9@3540_g N_VDD_Mp9@3540_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3539 N_OUT9_Mn9@3539_d N_OUT8_Mn9@3539_g N_VSS_Mn9@3539_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3538 N_OUT9_Mn9@3538_d N_OUT8_Mn9@3538_g N_VSS_Mn9@3538_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3539 N_OUT9_Mp9@3539_d N_OUT8_Mp9@3539_g N_VDD_Mp9@3539_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3538 N_OUT9_Mp9@3538_d N_OUT8_Mp9@3538_g N_VDD_Mp9@3538_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3537 N_OUT9_Mn9@3537_d N_OUT8_Mn9@3537_g N_VSS_Mn9@3537_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3536 N_OUT9_Mn9@3536_d N_OUT8_Mn9@3536_g N_VSS_Mn9@3536_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3537 N_OUT9_Mp9@3537_d N_OUT8_Mp9@3537_g N_VDD_Mp9@3537_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3536 N_OUT9_Mp9@3536_d N_OUT8_Mp9@3536_g N_VDD_Mp9@3536_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3535 N_OUT9_Mn9@3535_d N_OUT8_Mn9@3535_g N_VSS_Mn9@3535_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3534 N_OUT9_Mn9@3534_d N_OUT8_Mn9@3534_g N_VSS_Mn9@3534_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3535 N_OUT9_Mp9@3535_d N_OUT8_Mp9@3535_g N_VDD_Mp9@3535_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3534 N_OUT9_Mp9@3534_d N_OUT8_Mp9@3534_g N_VDD_Mp9@3534_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3533 N_OUT9_Mn9@3533_d N_OUT8_Mn9@3533_g N_VSS_Mn9@3533_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3532 N_OUT9_Mn9@3532_d N_OUT8_Mn9@3532_g N_VSS_Mn9@3532_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3533 N_OUT9_Mp9@3533_d N_OUT8_Mp9@3533_g N_VDD_Mp9@3533_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3532 N_OUT9_Mp9@3532_d N_OUT8_Mp9@3532_g N_VDD_Mp9@3532_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3531 N_OUT9_Mn9@3531_d N_OUT8_Mn9@3531_g N_VSS_Mn9@3531_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3530 N_OUT9_Mn9@3530_d N_OUT8_Mn9@3530_g N_VSS_Mn9@3530_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3531 N_OUT9_Mp9@3531_d N_OUT8_Mp9@3531_g N_VDD_Mp9@3531_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3530 N_OUT9_Mp9@3530_d N_OUT8_Mp9@3530_g N_VDD_Mp9@3530_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3529 N_OUT9_Mn9@3529_d N_OUT8_Mn9@3529_g N_VSS_Mn9@3529_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3528 N_OUT9_Mn9@3528_d N_OUT8_Mn9@3528_g N_VSS_Mn9@3528_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3529 N_OUT9_Mp9@3529_d N_OUT8_Mp9@3529_g N_VDD_Mp9@3529_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3528 N_OUT9_Mp9@3528_d N_OUT8_Mp9@3528_g N_VDD_Mp9@3528_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3527 N_OUT9_Mn9@3527_d N_OUT8_Mn9@3527_g N_VSS_Mn9@3527_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3526 N_OUT9_Mn9@3526_d N_OUT8_Mn9@3526_g N_VSS_Mn9@3526_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3527 N_OUT9_Mp9@3527_d N_OUT8_Mp9@3527_g N_VDD_Mp9@3527_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3526 N_OUT9_Mp9@3526_d N_OUT8_Mp9@3526_g N_VDD_Mp9@3526_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3525 N_OUT9_Mn9@3525_d N_OUT8_Mn9@3525_g N_VSS_Mn9@3525_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3524 N_OUT9_Mn9@3524_d N_OUT8_Mn9@3524_g N_VSS_Mn9@3524_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3525 N_OUT9_Mp9@3525_d N_OUT8_Mp9@3525_g N_VDD_Mp9@3525_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3524 N_OUT9_Mp9@3524_d N_OUT8_Mp9@3524_g N_VDD_Mp9@3524_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3523 N_OUT9_Mn9@3523_d N_OUT8_Mn9@3523_g N_VSS_Mn9@3523_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3522 N_OUT9_Mn9@3522_d N_OUT8_Mn9@3522_g N_VSS_Mn9@3522_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3523 N_OUT9_Mp9@3523_d N_OUT8_Mp9@3523_g N_VDD_Mp9@3523_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3522 N_OUT9_Mp9@3522_d N_OUT8_Mp9@3522_g N_VDD_Mp9@3522_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3521 N_OUT9_Mn9@3521_d N_OUT8_Mn9@3521_g N_VSS_Mn9@3521_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3520 N_OUT9_Mn9@3520_d N_OUT8_Mn9@3520_g N_VSS_Mn9@3520_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3521 N_OUT9_Mp9@3521_d N_OUT8_Mp9@3521_g N_VDD_Mp9@3521_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3520 N_OUT9_Mp9@3520_d N_OUT8_Mp9@3520_g N_VDD_Mp9@3520_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3519 N_OUT9_Mn9@3519_d N_OUT8_Mn9@3519_g N_VSS_Mn9@3519_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3518 N_OUT9_Mn9@3518_d N_OUT8_Mn9@3518_g N_VSS_Mn9@3518_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3519 N_OUT9_Mp9@3519_d N_OUT8_Mp9@3519_g N_VDD_Mp9@3519_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3518 N_OUT9_Mp9@3518_d N_OUT8_Mp9@3518_g N_VDD_Mp9@3518_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3517 N_OUT9_Mn9@3517_d N_OUT8_Mn9@3517_g N_VSS_Mn9@3517_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3516 N_OUT9_Mn9@3516_d N_OUT8_Mn9@3516_g N_VSS_Mn9@3516_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3517 N_OUT9_Mp9@3517_d N_OUT8_Mp9@3517_g N_VDD_Mp9@3517_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3516 N_OUT9_Mp9@3516_d N_OUT8_Mp9@3516_g N_VDD_Mp9@3516_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3515 N_OUT9_Mn9@3515_d N_OUT8_Mn9@3515_g N_VSS_Mn9@3515_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3514 N_OUT9_Mn9@3514_d N_OUT8_Mn9@3514_g N_VSS_Mn9@3514_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3515 N_OUT9_Mp9@3515_d N_OUT8_Mp9@3515_g N_VDD_Mp9@3515_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3514 N_OUT9_Mp9@3514_d N_OUT8_Mp9@3514_g N_VDD_Mp9@3514_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3513 N_OUT9_Mn9@3513_d N_OUT8_Mn9@3513_g N_VSS_Mn9@3513_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3512 N_OUT9_Mn9@3512_d N_OUT8_Mn9@3512_g N_VSS_Mn9@3512_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3513 N_OUT9_Mp9@3513_d N_OUT8_Mp9@3513_g N_VDD_Mp9@3513_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3512 N_OUT9_Mp9@3512_d N_OUT8_Mp9@3512_g N_VDD_Mp9@3512_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3511 N_OUT9_Mn9@3511_d N_OUT8_Mn9@3511_g N_VSS_Mn9@3511_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3510 N_OUT9_Mn9@3510_d N_OUT8_Mn9@3510_g N_VSS_Mn9@3510_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3511 N_OUT9_Mp9@3511_d N_OUT8_Mp9@3511_g N_VDD_Mp9@3511_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3510 N_OUT9_Mp9@3510_d N_OUT8_Mp9@3510_g N_VDD_Mp9@3510_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3509 N_OUT9_Mn9@3509_d N_OUT8_Mn9@3509_g N_VSS_Mn9@3509_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3508 N_OUT9_Mn9@3508_d N_OUT8_Mn9@3508_g N_VSS_Mn9@3508_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3509 N_OUT9_Mp9@3509_d N_OUT8_Mp9@3509_g N_VDD_Mp9@3509_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3508 N_OUT9_Mp9@3508_d N_OUT8_Mp9@3508_g N_VDD_Mp9@3508_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3507 N_OUT9_Mn9@3507_d N_OUT8_Mn9@3507_g N_VSS_Mn9@3507_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3506 N_OUT9_Mn9@3506_d N_OUT8_Mn9@3506_g N_VSS_Mn9@3506_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3507 N_OUT9_Mp9@3507_d N_OUT8_Mp9@3507_g N_VDD_Mp9@3507_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3506 N_OUT9_Mp9@3506_d N_OUT8_Mp9@3506_g N_VDD_Mp9@3506_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3505 N_OUT9_Mn9@3505_d N_OUT8_Mn9@3505_g N_VSS_Mn9@3505_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3504 N_OUT9_Mn9@3504_d N_OUT8_Mn9@3504_g N_VSS_Mn9@3504_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3505 N_OUT9_Mp9@3505_d N_OUT8_Mp9@3505_g N_VDD_Mp9@3505_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3504 N_OUT9_Mp9@3504_d N_OUT8_Mp9@3504_g N_VDD_Mp9@3504_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3503 N_OUT9_Mn9@3503_d N_OUT8_Mn9@3503_g N_VSS_Mn9@3503_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3502 N_OUT9_Mn9@3502_d N_OUT8_Mn9@3502_g N_VSS_Mn9@3502_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3503 N_OUT9_Mp9@3503_d N_OUT8_Mp9@3503_g N_VDD_Mp9@3503_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3502 N_OUT9_Mp9@3502_d N_OUT8_Mp9@3502_g N_VDD_Mp9@3502_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3501 N_OUT9_Mn9@3501_d N_OUT8_Mn9@3501_g N_VSS_Mn9@3501_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3500 N_OUT9_Mn9@3500_d N_OUT8_Mn9@3500_g N_VSS_Mn9@3500_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3501 N_OUT9_Mp9@3501_d N_OUT8_Mp9@3501_g N_VDD_Mp9@3501_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3500 N_OUT9_Mp9@3500_d N_OUT8_Mp9@3500_g N_VDD_Mp9@3500_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3499 N_OUT9_Mn9@3499_d N_OUT8_Mn9@3499_g N_VSS_Mn9@3499_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3498 N_OUT9_Mn9@3498_d N_OUT8_Mn9@3498_g N_VSS_Mn9@3498_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3499 N_OUT9_Mp9@3499_d N_OUT8_Mp9@3499_g N_VDD_Mp9@3499_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3498 N_OUT9_Mp9@3498_d N_OUT8_Mp9@3498_g N_VDD_Mp9@3498_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3497 N_OUT9_Mn9@3497_d N_OUT8_Mn9@3497_g N_VSS_Mn9@3497_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3496 N_OUT9_Mn9@3496_d N_OUT8_Mn9@3496_g N_VSS_Mn9@3496_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3497 N_OUT9_Mp9@3497_d N_OUT8_Mp9@3497_g N_VDD_Mp9@3497_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3496 N_OUT9_Mp9@3496_d N_OUT8_Mp9@3496_g N_VDD_Mp9@3496_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3495 N_OUT9_Mn9@3495_d N_OUT8_Mn9@3495_g N_VSS_Mn9@3495_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3494 N_OUT9_Mn9@3494_d N_OUT8_Mn9@3494_g N_VSS_Mn9@3494_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3495 N_OUT9_Mp9@3495_d N_OUT8_Mp9@3495_g N_VDD_Mp9@3495_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3494 N_OUT9_Mp9@3494_d N_OUT8_Mp9@3494_g N_VDD_Mp9@3494_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3493 N_OUT9_Mn9@3493_d N_OUT8_Mn9@3493_g N_VSS_Mn9@3493_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3492 N_OUT9_Mn9@3492_d N_OUT8_Mn9@3492_g N_VSS_Mn9@3492_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3493 N_OUT9_Mp9@3493_d N_OUT8_Mp9@3493_g N_VDD_Mp9@3493_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3492 N_OUT9_Mp9@3492_d N_OUT8_Mp9@3492_g N_VDD_Mp9@3492_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3491 N_OUT9_Mn9@3491_d N_OUT8_Mn9@3491_g N_VSS_Mn9@3491_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3490 N_OUT9_Mn9@3490_d N_OUT8_Mn9@3490_g N_VSS_Mn9@3490_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3491 N_OUT9_Mp9@3491_d N_OUT8_Mp9@3491_g N_VDD_Mp9@3491_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3490 N_OUT9_Mp9@3490_d N_OUT8_Mp9@3490_g N_VDD_Mp9@3490_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3489 N_OUT9_Mn9@3489_d N_OUT8_Mn9@3489_g N_VSS_Mn9@3489_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3488 N_OUT9_Mn9@3488_d N_OUT8_Mn9@3488_g N_VSS_Mn9@3488_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3489 N_OUT9_Mp9@3489_d N_OUT8_Mp9@3489_g N_VDD_Mp9@3489_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3488 N_OUT9_Mp9@3488_d N_OUT8_Mp9@3488_g N_VDD_Mp9@3488_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3487 N_OUT9_Mn9@3487_d N_OUT8_Mn9@3487_g N_VSS_Mn9@3487_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3486 N_OUT9_Mn9@3486_d N_OUT8_Mn9@3486_g N_VSS_Mn9@3486_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3487 N_OUT9_Mp9@3487_d N_OUT8_Mp9@3487_g N_VDD_Mp9@3487_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3486 N_OUT9_Mp9@3486_d N_OUT8_Mp9@3486_g N_VDD_Mp9@3486_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3485 N_OUT9_Mn9@3485_d N_OUT8_Mn9@3485_g N_VSS_Mn9@3485_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3484 N_OUT9_Mn9@3484_d N_OUT8_Mn9@3484_g N_VSS_Mn9@3484_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3485 N_OUT9_Mp9@3485_d N_OUT8_Mp9@3485_g N_VDD_Mp9@3485_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3484 N_OUT9_Mp9@3484_d N_OUT8_Mp9@3484_g N_VDD_Mp9@3484_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3483 N_OUT9_Mn9@3483_d N_OUT8_Mn9@3483_g N_VSS_Mn9@3483_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3482 N_OUT9_Mn9@3482_d N_OUT8_Mn9@3482_g N_VSS_Mn9@3482_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3483 N_OUT9_Mp9@3483_d N_OUT8_Mp9@3483_g N_VDD_Mp9@3483_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3482 N_OUT9_Mp9@3482_d N_OUT8_Mp9@3482_g N_VDD_Mp9@3482_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3481 N_OUT9_Mn9@3481_d N_OUT8_Mn9@3481_g N_VSS_Mn9@3481_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3480 N_OUT9_Mn9@3480_d N_OUT8_Mn9@3480_g N_VSS_Mn9@3480_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3481 N_OUT9_Mp9@3481_d N_OUT8_Mp9@3481_g N_VDD_Mp9@3481_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3480 N_OUT9_Mp9@3480_d N_OUT8_Mp9@3480_g N_VDD_Mp9@3480_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3479 N_OUT9_Mn9@3479_d N_OUT8_Mn9@3479_g N_VSS_Mn9@3479_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3478 N_OUT9_Mn9@3478_d N_OUT8_Mn9@3478_g N_VSS_Mn9@3478_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3479 N_OUT9_Mp9@3479_d N_OUT8_Mp9@3479_g N_VDD_Mp9@3479_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3478 N_OUT9_Mp9@3478_d N_OUT8_Mp9@3478_g N_VDD_Mp9@3478_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3477 N_OUT9_Mn9@3477_d N_OUT8_Mn9@3477_g N_VSS_Mn9@3477_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3476 N_OUT9_Mn9@3476_d N_OUT8_Mn9@3476_g N_VSS_Mn9@3476_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3477 N_OUT9_Mp9@3477_d N_OUT8_Mp9@3477_g N_VDD_Mp9@3477_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3476 N_OUT9_Mp9@3476_d N_OUT8_Mp9@3476_g N_VDD_Mp9@3476_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3475 N_OUT9_Mn9@3475_d N_OUT8_Mn9@3475_g N_VSS_Mn9@3475_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3474 N_OUT9_Mn9@3474_d N_OUT8_Mn9@3474_g N_VSS_Mn9@3474_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3475 N_OUT9_Mp9@3475_d N_OUT8_Mp9@3475_g N_VDD_Mp9@3475_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3474 N_OUT9_Mp9@3474_d N_OUT8_Mp9@3474_g N_VDD_Mp9@3474_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3473 N_OUT9_Mn9@3473_d N_OUT8_Mn9@3473_g N_VSS_Mn9@3473_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3472 N_OUT9_Mn9@3472_d N_OUT8_Mn9@3472_g N_VSS_Mn9@3472_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3473 N_OUT9_Mp9@3473_d N_OUT8_Mp9@3473_g N_VDD_Mp9@3473_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3472 N_OUT9_Mp9@3472_d N_OUT8_Mp9@3472_g N_VDD_Mp9@3472_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3471 N_OUT9_Mn9@3471_d N_OUT8_Mn9@3471_g N_VSS_Mn9@3471_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3470 N_OUT9_Mn9@3470_d N_OUT8_Mn9@3470_g N_VSS_Mn9@3470_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3471 N_OUT9_Mp9@3471_d N_OUT8_Mp9@3471_g N_VDD_Mp9@3471_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3470 N_OUT9_Mp9@3470_d N_OUT8_Mp9@3470_g N_VDD_Mp9@3470_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3469 N_OUT9_Mn9@3469_d N_OUT8_Mn9@3469_g N_VSS_Mn9@3469_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3468 N_OUT9_Mn9@3468_d N_OUT8_Mn9@3468_g N_VSS_Mn9@3468_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3469 N_OUT9_Mp9@3469_d N_OUT8_Mp9@3469_g N_VDD_Mp9@3469_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3468 N_OUT9_Mp9@3468_d N_OUT8_Mp9@3468_g N_VDD_Mp9@3468_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3467 N_OUT9_Mn9@3467_d N_OUT8_Mn9@3467_g N_VSS_Mn9@3467_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3466 N_OUT9_Mn9@3466_d N_OUT8_Mn9@3466_g N_VSS_Mn9@3466_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3467 N_OUT9_Mp9@3467_d N_OUT8_Mp9@3467_g N_VDD_Mp9@3467_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3466 N_OUT9_Mp9@3466_d N_OUT8_Mp9@3466_g N_VDD_Mp9@3466_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3465 N_OUT9_Mn9@3465_d N_OUT8_Mn9@3465_g N_VSS_Mn9@3465_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3464 N_OUT9_Mn9@3464_d N_OUT8_Mn9@3464_g N_VSS_Mn9@3464_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3465 N_OUT9_Mp9@3465_d N_OUT8_Mp9@3465_g N_VDD_Mp9@3465_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3464 N_OUT9_Mp9@3464_d N_OUT8_Mp9@3464_g N_VDD_Mp9@3464_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3463 N_OUT9_Mn9@3463_d N_OUT8_Mn9@3463_g N_VSS_Mn9@3463_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3462 N_OUT9_Mn9@3462_d N_OUT8_Mn9@3462_g N_VSS_Mn9@3462_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3463 N_OUT9_Mp9@3463_d N_OUT8_Mp9@3463_g N_VDD_Mp9@3463_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3462 N_OUT9_Mp9@3462_d N_OUT8_Mp9@3462_g N_VDD_Mp9@3462_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3461 N_OUT9_Mn9@3461_d N_OUT8_Mn9@3461_g N_VSS_Mn9@3461_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3460 N_OUT9_Mn9@3460_d N_OUT8_Mn9@3460_g N_VSS_Mn9@3460_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3461 N_OUT9_Mp9@3461_d N_OUT8_Mp9@3461_g N_VDD_Mp9@3461_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3460 N_OUT9_Mp9@3460_d N_OUT8_Mp9@3460_g N_VDD_Mp9@3460_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3459 N_OUT9_Mn9@3459_d N_OUT8_Mn9@3459_g N_VSS_Mn9@3459_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3458 N_OUT9_Mn9@3458_d N_OUT8_Mn9@3458_g N_VSS_Mn9@3458_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3459 N_OUT9_Mp9@3459_d N_OUT8_Mp9@3459_g N_VDD_Mp9@3459_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3458 N_OUT9_Mp9@3458_d N_OUT8_Mp9@3458_g N_VDD_Mp9@3458_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3457 N_OUT9_Mn9@3457_d N_OUT8_Mn9@3457_g N_VSS_Mn9@3457_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3456 N_OUT9_Mn9@3456_d N_OUT8_Mn9@3456_g N_VSS_Mn9@3456_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3457 N_OUT9_Mp9@3457_d N_OUT8_Mp9@3457_g N_VDD_Mp9@3457_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3456 N_OUT9_Mp9@3456_d N_OUT8_Mp9@3456_g N_VDD_Mp9@3456_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3455 N_OUT9_Mn9@3455_d N_OUT8_Mn9@3455_g N_VSS_Mn9@3455_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3454 N_OUT9_Mn9@3454_d N_OUT8_Mn9@3454_g N_VSS_Mn9@3454_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3455 N_OUT9_Mp9@3455_d N_OUT8_Mp9@3455_g N_VDD_Mp9@3455_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3454 N_OUT9_Mp9@3454_d N_OUT8_Mp9@3454_g N_VDD_Mp9@3454_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3453 N_OUT9_Mn9@3453_d N_OUT8_Mn9@3453_g N_VSS_Mn9@3453_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3452 N_OUT9_Mn9@3452_d N_OUT8_Mn9@3452_g N_VSS_Mn9@3452_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3453 N_OUT9_Mp9@3453_d N_OUT8_Mp9@3453_g N_VDD_Mp9@3453_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3452 N_OUT9_Mp9@3452_d N_OUT8_Mp9@3452_g N_VDD_Mp9@3452_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3451 N_OUT9_Mn9@3451_d N_OUT8_Mn9@3451_g N_VSS_Mn9@3451_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3450 N_OUT9_Mn9@3450_d N_OUT8_Mn9@3450_g N_VSS_Mn9@3450_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3451 N_OUT9_Mp9@3451_d N_OUT8_Mp9@3451_g N_VDD_Mp9@3451_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3450 N_OUT9_Mp9@3450_d N_OUT8_Mp9@3450_g N_VDD_Mp9@3450_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3449 N_OUT9_Mn9@3449_d N_OUT8_Mn9@3449_g N_VSS_Mn9@3449_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3448 N_OUT9_Mn9@3448_d N_OUT8_Mn9@3448_g N_VSS_Mn9@3448_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3449 N_OUT9_Mp9@3449_d N_OUT8_Mp9@3449_g N_VDD_Mp9@3449_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3448 N_OUT9_Mp9@3448_d N_OUT8_Mp9@3448_g N_VDD_Mp9@3448_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3447 N_OUT9_Mn9@3447_d N_OUT8_Mn9@3447_g N_VSS_Mn9@3447_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3446 N_OUT9_Mn9@3446_d N_OUT8_Mn9@3446_g N_VSS_Mn9@3446_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3447 N_OUT9_Mp9@3447_d N_OUT8_Mp9@3447_g N_VDD_Mp9@3447_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3446 N_OUT9_Mp9@3446_d N_OUT8_Mp9@3446_g N_VDD_Mp9@3446_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3445 N_OUT9_Mn9@3445_d N_OUT8_Mn9@3445_g N_VSS_Mn9@3445_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3444 N_OUT9_Mn9@3444_d N_OUT8_Mn9@3444_g N_VSS_Mn9@3444_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3445 N_OUT9_Mp9@3445_d N_OUT8_Mp9@3445_g N_VDD_Mp9@3445_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3444 N_OUT9_Mp9@3444_d N_OUT8_Mp9@3444_g N_VDD_Mp9@3444_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3443 N_OUT9_Mn9@3443_d N_OUT8_Mn9@3443_g N_VSS_Mn9@3443_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3442 N_OUT9_Mn9@3442_d N_OUT8_Mn9@3442_g N_VSS_Mn9@3442_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3443 N_OUT9_Mp9@3443_d N_OUT8_Mp9@3443_g N_VDD_Mp9@3443_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3442 N_OUT9_Mp9@3442_d N_OUT8_Mp9@3442_g N_VDD_Mp9@3442_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3441 N_OUT9_Mn9@3441_d N_OUT8_Mn9@3441_g N_VSS_Mn9@3441_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3440 N_OUT9_Mn9@3440_d N_OUT8_Mn9@3440_g N_VSS_Mn9@3440_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3441 N_OUT9_Mp9@3441_d N_OUT8_Mp9@3441_g N_VDD_Mp9@3441_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3440 N_OUT9_Mp9@3440_d N_OUT8_Mp9@3440_g N_VDD_Mp9@3440_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3439 N_OUT9_Mn9@3439_d N_OUT8_Mn9@3439_g N_VSS_Mn9@3439_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3438 N_OUT9_Mn9@3438_d N_OUT8_Mn9@3438_g N_VSS_Mn9@3438_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3439 N_OUT9_Mp9@3439_d N_OUT8_Mp9@3439_g N_VDD_Mp9@3439_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3438 N_OUT9_Mp9@3438_d N_OUT8_Mp9@3438_g N_VDD_Mp9@3438_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3437 N_OUT9_Mn9@3437_d N_OUT8_Mn9@3437_g N_VSS_Mn9@3437_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3436 N_OUT9_Mn9@3436_d N_OUT8_Mn9@3436_g N_VSS_Mn9@3436_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3437 N_OUT9_Mp9@3437_d N_OUT8_Mp9@3437_g N_VDD_Mp9@3437_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3436 N_OUT9_Mp9@3436_d N_OUT8_Mp9@3436_g N_VDD_Mp9@3436_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3435 N_OUT9_Mn9@3435_d N_OUT8_Mn9@3435_g N_VSS_Mn9@3435_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3434 N_OUT9_Mn9@3434_d N_OUT8_Mn9@3434_g N_VSS_Mn9@3434_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3435 N_OUT9_Mp9@3435_d N_OUT8_Mp9@3435_g N_VDD_Mp9@3435_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3434 N_OUT9_Mp9@3434_d N_OUT8_Mp9@3434_g N_VDD_Mp9@3434_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3433 N_OUT9_Mn9@3433_d N_OUT8_Mn9@3433_g N_VSS_Mn9@3433_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3432 N_OUT9_Mn9@3432_d N_OUT8_Mn9@3432_g N_VSS_Mn9@3432_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3433 N_OUT9_Mp9@3433_d N_OUT8_Mp9@3433_g N_VDD_Mp9@3433_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3432 N_OUT9_Mp9@3432_d N_OUT8_Mp9@3432_g N_VDD_Mp9@3432_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3431 N_OUT9_Mn9@3431_d N_OUT8_Mn9@3431_g N_VSS_Mn9@3431_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3430 N_OUT9_Mn9@3430_d N_OUT8_Mn9@3430_g N_VSS_Mn9@3430_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3431 N_OUT9_Mp9@3431_d N_OUT8_Mp9@3431_g N_VDD_Mp9@3431_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3430 N_OUT9_Mp9@3430_d N_OUT8_Mp9@3430_g N_VDD_Mp9@3430_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3429 N_OUT9_Mn9@3429_d N_OUT8_Mn9@3429_g N_VSS_Mn9@3429_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3428 N_OUT9_Mn9@3428_d N_OUT8_Mn9@3428_g N_VSS_Mn9@3428_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3429 N_OUT9_Mp9@3429_d N_OUT8_Mp9@3429_g N_VDD_Mp9@3429_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3428 N_OUT9_Mp9@3428_d N_OUT8_Mp9@3428_g N_VDD_Mp9@3428_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3427 N_OUT9_Mn9@3427_d N_OUT8_Mn9@3427_g N_VSS_Mn9@3427_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3426 N_OUT9_Mn9@3426_d N_OUT8_Mn9@3426_g N_VSS_Mn9@3426_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3427 N_OUT9_Mp9@3427_d N_OUT8_Mp9@3427_g N_VDD_Mp9@3427_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3426 N_OUT9_Mp9@3426_d N_OUT8_Mp9@3426_g N_VDD_Mp9@3426_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3425 N_OUT9_Mn9@3425_d N_OUT8_Mn9@3425_g N_VSS_Mn9@3425_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3424 N_OUT9_Mn9@3424_d N_OUT8_Mn9@3424_g N_VSS_Mn9@3424_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3425 N_OUT9_Mp9@3425_d N_OUT8_Mp9@3425_g N_VDD_Mp9@3425_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3424 N_OUT9_Mp9@3424_d N_OUT8_Mp9@3424_g N_VDD_Mp9@3424_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3423 N_OUT9_Mn9@3423_d N_OUT8_Mn9@3423_g N_VSS_Mn9@3423_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3422 N_OUT9_Mn9@3422_d N_OUT8_Mn9@3422_g N_VSS_Mn9@3422_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3423 N_OUT9_Mp9@3423_d N_OUT8_Mp9@3423_g N_VDD_Mp9@3423_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3422 N_OUT9_Mp9@3422_d N_OUT8_Mp9@3422_g N_VDD_Mp9@3422_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3421 N_OUT9_Mn9@3421_d N_OUT8_Mn9@3421_g N_VSS_Mn9@3421_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3420 N_OUT9_Mn9@3420_d N_OUT8_Mn9@3420_g N_VSS_Mn9@3420_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3421 N_OUT9_Mp9@3421_d N_OUT8_Mp9@3421_g N_VDD_Mp9@3421_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3420 N_OUT9_Mp9@3420_d N_OUT8_Mp9@3420_g N_VDD_Mp9@3420_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3419 N_OUT9_Mn9@3419_d N_OUT8_Mn9@3419_g N_VSS_Mn9@3419_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3418 N_OUT9_Mn9@3418_d N_OUT8_Mn9@3418_g N_VSS_Mn9@3418_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3419 N_OUT9_Mp9@3419_d N_OUT8_Mp9@3419_g N_VDD_Mp9@3419_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3418 N_OUT9_Mp9@3418_d N_OUT8_Mp9@3418_g N_VDD_Mp9@3418_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3417 N_OUT9_Mn9@3417_d N_OUT8_Mn9@3417_g N_VSS_Mn9@3417_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3416 N_OUT9_Mn9@3416_d N_OUT8_Mn9@3416_g N_VSS_Mn9@3416_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3417 N_OUT9_Mp9@3417_d N_OUT8_Mp9@3417_g N_VDD_Mp9@3417_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3416 N_OUT9_Mp9@3416_d N_OUT8_Mp9@3416_g N_VDD_Mp9@3416_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3415 N_OUT9_Mn9@3415_d N_OUT8_Mn9@3415_g N_VSS_Mn9@3415_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3414 N_OUT9_Mn9@3414_d N_OUT8_Mn9@3414_g N_VSS_Mn9@3414_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3415 N_OUT9_Mp9@3415_d N_OUT8_Mp9@3415_g N_VDD_Mp9@3415_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3414 N_OUT9_Mp9@3414_d N_OUT8_Mp9@3414_g N_VDD_Mp9@3414_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3413 N_OUT9_Mn9@3413_d N_OUT8_Mn9@3413_g N_VSS_Mn9@3413_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3412 N_OUT9_Mn9@3412_d N_OUT8_Mn9@3412_g N_VSS_Mn9@3412_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3413 N_OUT9_Mp9@3413_d N_OUT8_Mp9@3413_g N_VDD_Mp9@3413_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3412 N_OUT9_Mp9@3412_d N_OUT8_Mp9@3412_g N_VDD_Mp9@3412_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3411 N_OUT9_Mn9@3411_d N_OUT8_Mn9@3411_g N_VSS_Mn9@3411_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3410 N_OUT9_Mn9@3410_d N_OUT8_Mn9@3410_g N_VSS_Mn9@3410_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3411 N_OUT9_Mp9@3411_d N_OUT8_Mp9@3411_g N_VDD_Mp9@3411_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3410 N_OUT9_Mp9@3410_d N_OUT8_Mp9@3410_g N_VDD_Mp9@3410_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3409 N_OUT9_Mn9@3409_d N_OUT8_Mn9@3409_g N_VSS_Mn9@3409_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3408 N_OUT9_Mn9@3408_d N_OUT8_Mn9@3408_g N_VSS_Mn9@3408_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3409 N_OUT9_Mp9@3409_d N_OUT8_Mp9@3409_g N_VDD_Mp9@3409_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3408 N_OUT9_Mp9@3408_d N_OUT8_Mp9@3408_g N_VDD_Mp9@3408_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3407 N_OUT9_Mn9@3407_d N_OUT8_Mn9@3407_g N_VSS_Mn9@3407_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3406 N_OUT9_Mn9@3406_d N_OUT8_Mn9@3406_g N_VSS_Mn9@3406_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3407 N_OUT9_Mp9@3407_d N_OUT8_Mp9@3407_g N_VDD_Mp9@3407_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3406 N_OUT9_Mp9@3406_d N_OUT8_Mp9@3406_g N_VDD_Mp9@3406_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3405 N_OUT9_Mn9@3405_d N_OUT8_Mn9@3405_g N_VSS_Mn9@3405_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3404 N_OUT9_Mn9@3404_d N_OUT8_Mn9@3404_g N_VSS_Mn9@3404_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3405 N_OUT9_Mp9@3405_d N_OUT8_Mp9@3405_g N_VDD_Mp9@3405_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3404 N_OUT9_Mp9@3404_d N_OUT8_Mp9@3404_g N_VDD_Mp9@3404_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3403 N_OUT9_Mn9@3403_d N_OUT8_Mn9@3403_g N_VSS_Mn9@3403_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3402 N_OUT9_Mn9@3402_d N_OUT8_Mn9@3402_g N_VSS_Mn9@3402_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3403 N_OUT9_Mp9@3403_d N_OUT8_Mp9@3403_g N_VDD_Mp9@3403_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3402 N_OUT9_Mp9@3402_d N_OUT8_Mp9@3402_g N_VDD_Mp9@3402_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3401 N_OUT9_Mn9@3401_d N_OUT8_Mn9@3401_g N_VSS_Mn9@3401_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3400 N_OUT9_Mn9@3400_d N_OUT8_Mn9@3400_g N_VSS_Mn9@3400_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3401 N_OUT9_Mp9@3401_d N_OUT8_Mp9@3401_g N_VDD_Mp9@3401_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3400 N_OUT9_Mp9@3400_d N_OUT8_Mp9@3400_g N_VDD_Mp9@3400_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3399 N_OUT9_Mn9@3399_d N_OUT8_Mn9@3399_g N_VSS_Mn9@3399_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3398 N_OUT9_Mn9@3398_d N_OUT8_Mn9@3398_g N_VSS_Mn9@3398_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3399 N_OUT9_Mp9@3399_d N_OUT8_Mp9@3399_g N_VDD_Mp9@3399_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3398 N_OUT9_Mp9@3398_d N_OUT8_Mp9@3398_g N_VDD_Mp9@3398_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3397 N_OUT9_Mn9@3397_d N_OUT8_Mn9@3397_g N_VSS_Mn9@3397_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3396 N_OUT9_Mn9@3396_d N_OUT8_Mn9@3396_g N_VSS_Mn9@3396_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3397 N_OUT9_Mp9@3397_d N_OUT8_Mp9@3397_g N_VDD_Mp9@3397_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3396 N_OUT9_Mp9@3396_d N_OUT8_Mp9@3396_g N_VDD_Mp9@3396_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3395 N_OUT9_Mn9@3395_d N_OUT8_Mn9@3395_g N_VSS_Mn9@3395_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3394 N_OUT9_Mn9@3394_d N_OUT8_Mn9@3394_g N_VSS_Mn9@3394_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3395 N_OUT9_Mp9@3395_d N_OUT8_Mp9@3395_g N_VDD_Mp9@3395_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3394 N_OUT9_Mp9@3394_d N_OUT8_Mp9@3394_g N_VDD_Mp9@3394_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3393 N_OUT9_Mn9@3393_d N_OUT8_Mn9@3393_g N_VSS_Mn9@3393_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3392 N_OUT9_Mn9@3392_d N_OUT8_Mn9@3392_g N_VSS_Mn9@3392_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3393 N_OUT9_Mp9@3393_d N_OUT8_Mp9@3393_g N_VDD_Mp9@3393_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3392 N_OUT9_Mp9@3392_d N_OUT8_Mp9@3392_g N_VDD_Mp9@3392_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3391 N_OUT9_Mn9@3391_d N_OUT8_Mn9@3391_g N_VSS_Mn9@3391_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3390 N_OUT9_Mn9@3390_d N_OUT8_Mn9@3390_g N_VSS_Mn9@3390_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3391 N_OUT9_Mp9@3391_d N_OUT8_Mp9@3391_g N_VDD_Mp9@3391_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3390 N_OUT9_Mp9@3390_d N_OUT8_Mp9@3390_g N_VDD_Mp9@3390_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3389 N_OUT9_Mn9@3389_d N_OUT8_Mn9@3389_g N_VSS_Mn9@3389_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3388 N_OUT9_Mn9@3388_d N_OUT8_Mn9@3388_g N_VSS_Mn9@3388_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3389 N_OUT9_Mp9@3389_d N_OUT8_Mp9@3389_g N_VDD_Mp9@3389_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3388 N_OUT9_Mp9@3388_d N_OUT8_Mp9@3388_g N_VDD_Mp9@3388_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3387 N_OUT9_Mn9@3387_d N_OUT8_Mn9@3387_g N_VSS_Mn9@3387_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3386 N_OUT9_Mn9@3386_d N_OUT8_Mn9@3386_g N_VSS_Mn9@3386_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3387 N_OUT9_Mp9@3387_d N_OUT8_Mp9@3387_g N_VDD_Mp9@3387_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3386 N_OUT9_Mp9@3386_d N_OUT8_Mp9@3386_g N_VDD_Mp9@3386_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3385 N_OUT9_Mn9@3385_d N_OUT8_Mn9@3385_g N_VSS_Mn9@3385_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3384 N_OUT9_Mn9@3384_d N_OUT8_Mn9@3384_g N_VSS_Mn9@3384_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3385 N_OUT9_Mp9@3385_d N_OUT8_Mp9@3385_g N_VDD_Mp9@3385_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3384 N_OUT9_Mp9@3384_d N_OUT8_Mp9@3384_g N_VDD_Mp9@3384_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3383 N_OUT9_Mn9@3383_d N_OUT8_Mn9@3383_g N_VSS_Mn9@3383_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3382 N_OUT9_Mn9@3382_d N_OUT8_Mn9@3382_g N_VSS_Mn9@3382_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3383 N_OUT9_Mp9@3383_d N_OUT8_Mp9@3383_g N_VDD_Mp9@3383_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3382 N_OUT9_Mp9@3382_d N_OUT8_Mp9@3382_g N_VDD_Mp9@3382_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3381 N_OUT9_Mn9@3381_d N_OUT8_Mn9@3381_g N_VSS_Mn9@3381_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3380 N_OUT9_Mn9@3380_d N_OUT8_Mn9@3380_g N_VSS_Mn9@3380_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3381 N_OUT9_Mp9@3381_d N_OUT8_Mp9@3381_g N_VDD_Mp9@3381_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3380 N_OUT9_Mp9@3380_d N_OUT8_Mp9@3380_g N_VDD_Mp9@3380_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3379 N_OUT9_Mn9@3379_d N_OUT8_Mn9@3379_g N_VSS_Mn9@3379_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3378 N_OUT9_Mn9@3378_d N_OUT8_Mn9@3378_g N_VSS_Mn9@3378_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3379 N_OUT9_Mp9@3379_d N_OUT8_Mp9@3379_g N_VDD_Mp9@3379_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3378 N_OUT9_Mp9@3378_d N_OUT8_Mp9@3378_g N_VDD_Mp9@3378_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3377 N_OUT9_Mn9@3377_d N_OUT8_Mn9@3377_g N_VSS_Mn9@3377_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3376 N_OUT9_Mn9@3376_d N_OUT8_Mn9@3376_g N_VSS_Mn9@3376_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3377 N_OUT9_Mp9@3377_d N_OUT8_Mp9@3377_g N_VDD_Mp9@3377_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3376 N_OUT9_Mp9@3376_d N_OUT8_Mp9@3376_g N_VDD_Mp9@3376_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3375 N_OUT9_Mn9@3375_d N_OUT8_Mn9@3375_g N_VSS_Mn9@3375_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3374 N_OUT9_Mn9@3374_d N_OUT8_Mn9@3374_g N_VSS_Mn9@3374_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3375 N_OUT9_Mp9@3375_d N_OUT8_Mp9@3375_g N_VDD_Mp9@3375_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3374 N_OUT9_Mp9@3374_d N_OUT8_Mp9@3374_g N_VDD_Mp9@3374_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3373 N_OUT9_Mn9@3373_d N_OUT8_Mn9@3373_g N_VSS_Mn9@3373_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3372 N_OUT9_Mn9@3372_d N_OUT8_Mn9@3372_g N_VSS_Mn9@3372_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3373 N_OUT9_Mp9@3373_d N_OUT8_Mp9@3373_g N_VDD_Mp9@3373_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3372 N_OUT9_Mp9@3372_d N_OUT8_Mp9@3372_g N_VDD_Mp9@3372_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3371 N_OUT9_Mn9@3371_d N_OUT8_Mn9@3371_g N_VSS_Mn9@3371_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3370 N_OUT9_Mn9@3370_d N_OUT8_Mn9@3370_g N_VSS_Mn9@3370_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3371 N_OUT9_Mp9@3371_d N_OUT8_Mp9@3371_g N_VDD_Mp9@3371_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3370 N_OUT9_Mp9@3370_d N_OUT8_Mp9@3370_g N_VDD_Mp9@3370_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3369 N_OUT9_Mn9@3369_d N_OUT8_Mn9@3369_g N_VSS_Mn9@3369_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3368 N_OUT9_Mn9@3368_d N_OUT8_Mn9@3368_g N_VSS_Mn9@3368_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3369 N_OUT9_Mp9@3369_d N_OUT8_Mp9@3369_g N_VDD_Mp9@3369_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3368 N_OUT9_Mp9@3368_d N_OUT8_Mp9@3368_g N_VDD_Mp9@3368_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3367 N_OUT9_Mn9@3367_d N_OUT8_Mn9@3367_g N_VSS_Mn9@3367_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3366 N_OUT9_Mn9@3366_d N_OUT8_Mn9@3366_g N_VSS_Mn9@3366_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3367 N_OUT9_Mp9@3367_d N_OUT8_Mp9@3367_g N_VDD_Mp9@3367_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3366 N_OUT9_Mp9@3366_d N_OUT8_Mp9@3366_g N_VDD_Mp9@3366_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3365 N_OUT9_Mn9@3365_d N_OUT8_Mn9@3365_g N_VSS_Mn9@3365_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3364 N_OUT9_Mn9@3364_d N_OUT8_Mn9@3364_g N_VSS_Mn9@3364_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3365 N_OUT9_Mp9@3365_d N_OUT8_Mp9@3365_g N_VDD_Mp9@3365_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3364 N_OUT9_Mp9@3364_d N_OUT8_Mp9@3364_g N_VDD_Mp9@3364_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3363 N_OUT9_Mn9@3363_d N_OUT8_Mn9@3363_g N_VSS_Mn9@3363_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3362 N_OUT9_Mn9@3362_d N_OUT8_Mn9@3362_g N_VSS_Mn9@3362_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3363 N_OUT9_Mp9@3363_d N_OUT8_Mp9@3363_g N_VDD_Mp9@3363_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3362 N_OUT9_Mp9@3362_d N_OUT8_Mp9@3362_g N_VDD_Mp9@3362_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3361 N_OUT9_Mn9@3361_d N_OUT8_Mn9@3361_g N_VSS_Mn9@3361_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3360 N_OUT9_Mn9@3360_d N_OUT8_Mn9@3360_g N_VSS_Mn9@3360_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3361 N_OUT9_Mp9@3361_d N_OUT8_Mp9@3361_g N_VDD_Mp9@3361_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3360 N_OUT9_Mp9@3360_d N_OUT8_Mp9@3360_g N_VDD_Mp9@3360_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3359 N_OUT9_Mn9@3359_d N_OUT8_Mn9@3359_g N_VSS_Mn9@3359_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3358 N_OUT9_Mn9@3358_d N_OUT8_Mn9@3358_g N_VSS_Mn9@3358_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3359 N_OUT9_Mp9@3359_d N_OUT8_Mp9@3359_g N_VDD_Mp9@3359_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3358 N_OUT9_Mp9@3358_d N_OUT8_Mp9@3358_g N_VDD_Mp9@3358_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3357 N_OUT9_Mn9@3357_d N_OUT8_Mn9@3357_g N_VSS_Mn9@3357_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3356 N_OUT9_Mn9@3356_d N_OUT8_Mn9@3356_g N_VSS_Mn9@3356_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3357 N_OUT9_Mp9@3357_d N_OUT8_Mp9@3357_g N_VDD_Mp9@3357_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3356 N_OUT9_Mp9@3356_d N_OUT8_Mp9@3356_g N_VDD_Mp9@3356_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3355 N_OUT9_Mn9@3355_d N_OUT8_Mn9@3355_g N_VSS_Mn9@3355_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3354 N_OUT9_Mn9@3354_d N_OUT8_Mn9@3354_g N_VSS_Mn9@3354_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3355 N_OUT9_Mp9@3355_d N_OUT8_Mp9@3355_g N_VDD_Mp9@3355_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3354 N_OUT9_Mp9@3354_d N_OUT8_Mp9@3354_g N_VDD_Mp9@3354_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3353 N_OUT9_Mn9@3353_d N_OUT8_Mn9@3353_g N_VSS_Mn9@3353_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3352 N_OUT9_Mn9@3352_d N_OUT8_Mn9@3352_g N_VSS_Mn9@3352_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3353 N_OUT9_Mp9@3353_d N_OUT8_Mp9@3353_g N_VDD_Mp9@3353_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3352 N_OUT9_Mp9@3352_d N_OUT8_Mp9@3352_g N_VDD_Mp9@3352_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3351 N_OUT9_Mn9@3351_d N_OUT8_Mn9@3351_g N_VSS_Mn9@3351_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3350 N_OUT9_Mn9@3350_d N_OUT8_Mn9@3350_g N_VSS_Mn9@3350_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3351 N_OUT9_Mp9@3351_d N_OUT8_Mp9@3351_g N_VDD_Mp9@3351_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3350 N_OUT9_Mp9@3350_d N_OUT8_Mp9@3350_g N_VDD_Mp9@3350_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3349 N_OUT9_Mn9@3349_d N_OUT8_Mn9@3349_g N_VSS_Mn9@3349_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3348 N_OUT9_Mn9@3348_d N_OUT8_Mn9@3348_g N_VSS_Mn9@3348_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3349 N_OUT9_Mp9@3349_d N_OUT8_Mp9@3349_g N_VDD_Mp9@3349_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3348 N_OUT9_Mp9@3348_d N_OUT8_Mp9@3348_g N_VDD_Mp9@3348_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3347 N_OUT9_Mn9@3347_d N_OUT8_Mn9@3347_g N_VSS_Mn9@3347_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3346 N_OUT9_Mn9@3346_d N_OUT8_Mn9@3346_g N_VSS_Mn9@3346_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3347 N_OUT9_Mp9@3347_d N_OUT8_Mp9@3347_g N_VDD_Mp9@3347_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3346 N_OUT9_Mp9@3346_d N_OUT8_Mp9@3346_g N_VDD_Mp9@3346_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3345 N_OUT9_Mn9@3345_d N_OUT8_Mn9@3345_g N_VSS_Mn9@3345_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3344 N_OUT9_Mn9@3344_d N_OUT8_Mn9@3344_g N_VSS_Mn9@3344_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3345 N_OUT9_Mp9@3345_d N_OUT8_Mp9@3345_g N_VDD_Mp9@3345_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3344 N_OUT9_Mp9@3344_d N_OUT8_Mp9@3344_g N_VDD_Mp9@3344_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3343 N_OUT9_Mn9@3343_d N_OUT8_Mn9@3343_g N_VSS_Mn9@3343_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3342 N_OUT9_Mn9@3342_d N_OUT8_Mn9@3342_g N_VSS_Mn9@3342_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3343 N_OUT9_Mp9@3343_d N_OUT8_Mp9@3343_g N_VDD_Mp9@3343_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3342 N_OUT9_Mp9@3342_d N_OUT8_Mp9@3342_g N_VDD_Mp9@3342_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3341 N_OUT9_Mn9@3341_d N_OUT8_Mn9@3341_g N_VSS_Mn9@3341_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3340 N_OUT9_Mn9@3340_d N_OUT8_Mn9@3340_g N_VSS_Mn9@3340_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3341 N_OUT9_Mp9@3341_d N_OUT8_Mp9@3341_g N_VDD_Mp9@3341_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3340 N_OUT9_Mp9@3340_d N_OUT8_Mp9@3340_g N_VDD_Mp9@3340_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3339 N_OUT9_Mn9@3339_d N_OUT8_Mn9@3339_g N_VSS_Mn9@3339_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3338 N_OUT9_Mn9@3338_d N_OUT8_Mn9@3338_g N_VSS_Mn9@3338_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3339 N_OUT9_Mp9@3339_d N_OUT8_Mp9@3339_g N_VDD_Mp9@3339_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3338 N_OUT9_Mp9@3338_d N_OUT8_Mp9@3338_g N_VDD_Mp9@3338_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3337 N_OUT9_Mn9@3337_d N_OUT8_Mn9@3337_g N_VSS_Mn9@3337_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3336 N_OUT9_Mn9@3336_d N_OUT8_Mn9@3336_g N_VSS_Mn9@3336_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3337 N_OUT9_Mp9@3337_d N_OUT8_Mp9@3337_g N_VDD_Mp9@3337_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3336 N_OUT9_Mp9@3336_d N_OUT8_Mp9@3336_g N_VDD_Mp9@3336_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3335 N_OUT9_Mn9@3335_d N_OUT8_Mn9@3335_g N_VSS_Mn9@3335_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3334 N_OUT9_Mn9@3334_d N_OUT8_Mn9@3334_g N_VSS_Mn9@3334_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3335 N_OUT9_Mp9@3335_d N_OUT8_Mp9@3335_g N_VDD_Mp9@3335_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3334 N_OUT9_Mp9@3334_d N_OUT8_Mp9@3334_g N_VDD_Mp9@3334_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3333 N_OUT9_Mn9@3333_d N_OUT8_Mn9@3333_g N_VSS_Mn9@3333_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3332 N_OUT9_Mn9@3332_d N_OUT8_Mn9@3332_g N_VSS_Mn9@3332_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3333 N_OUT9_Mp9@3333_d N_OUT8_Mp9@3333_g N_VDD_Mp9@3333_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3332 N_OUT9_Mp9@3332_d N_OUT8_Mp9@3332_g N_VDD_Mp9@3332_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3331 N_OUT9_Mn9@3331_d N_OUT8_Mn9@3331_g N_VSS_Mn9@3331_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3330 N_OUT9_Mn9@3330_d N_OUT8_Mn9@3330_g N_VSS_Mn9@3330_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3331 N_OUT9_Mp9@3331_d N_OUT8_Mp9@3331_g N_VDD_Mp9@3331_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3330 N_OUT9_Mp9@3330_d N_OUT8_Mp9@3330_g N_VDD_Mp9@3330_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3329 N_OUT9_Mn9@3329_d N_OUT8_Mn9@3329_g N_VSS_Mn9@3329_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3328 N_OUT9_Mn9@3328_d N_OUT8_Mn9@3328_g N_VSS_Mn9@3328_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3329 N_OUT9_Mp9@3329_d N_OUT8_Mp9@3329_g N_VDD_Mp9@3329_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3328 N_OUT9_Mp9@3328_d N_OUT8_Mp9@3328_g N_VDD_Mp9@3328_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3327 N_OUT9_Mn9@3327_d N_OUT8_Mn9@3327_g N_VSS_Mn9@3327_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3326 N_OUT9_Mn9@3326_d N_OUT8_Mn9@3326_g N_VSS_Mn9@3326_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3327 N_OUT9_Mp9@3327_d N_OUT8_Mp9@3327_g N_VDD_Mp9@3327_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3326 N_OUT9_Mp9@3326_d N_OUT8_Mp9@3326_g N_VDD_Mp9@3326_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3325 N_OUT9_Mn9@3325_d N_OUT8_Mn9@3325_g N_VSS_Mn9@3325_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3324 N_OUT9_Mn9@3324_d N_OUT8_Mn9@3324_g N_VSS_Mn9@3324_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3325 N_OUT9_Mp9@3325_d N_OUT8_Mp9@3325_g N_VDD_Mp9@3325_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3324 N_OUT9_Mp9@3324_d N_OUT8_Mp9@3324_g N_VDD_Mp9@3324_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3323 N_OUT9_Mn9@3323_d N_OUT8_Mn9@3323_g N_VSS_Mn9@3323_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3322 N_OUT9_Mn9@3322_d N_OUT8_Mn9@3322_g N_VSS_Mn9@3322_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3323 N_OUT9_Mp9@3323_d N_OUT8_Mp9@3323_g N_VDD_Mp9@3323_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3322 N_OUT9_Mp9@3322_d N_OUT8_Mp9@3322_g N_VDD_Mp9@3322_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3321 N_OUT9_Mn9@3321_d N_OUT8_Mn9@3321_g N_VSS_Mn9@3321_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3320 N_OUT9_Mn9@3320_d N_OUT8_Mn9@3320_g N_VSS_Mn9@3320_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3321 N_OUT9_Mp9@3321_d N_OUT8_Mp9@3321_g N_VDD_Mp9@3321_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3320 N_OUT9_Mp9@3320_d N_OUT8_Mp9@3320_g N_VDD_Mp9@3320_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3319 N_OUT9_Mn9@3319_d N_OUT8_Mn9@3319_g N_VSS_Mn9@3319_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3318 N_OUT9_Mn9@3318_d N_OUT8_Mn9@3318_g N_VSS_Mn9@3318_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3319 N_OUT9_Mp9@3319_d N_OUT8_Mp9@3319_g N_VDD_Mp9@3319_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3318 N_OUT9_Mp9@3318_d N_OUT8_Mp9@3318_g N_VDD_Mp9@3318_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3317 N_OUT9_Mn9@3317_d N_OUT8_Mn9@3317_g N_VSS_Mn9@3317_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3316 N_OUT9_Mn9@3316_d N_OUT8_Mn9@3316_g N_VSS_Mn9@3316_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3317 N_OUT9_Mp9@3317_d N_OUT8_Mp9@3317_g N_VDD_Mp9@3317_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3316 N_OUT9_Mp9@3316_d N_OUT8_Mp9@3316_g N_VDD_Mp9@3316_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3315 N_OUT9_Mn9@3315_d N_OUT8_Mn9@3315_g N_VSS_Mn9@3315_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3314 N_OUT9_Mn9@3314_d N_OUT8_Mn9@3314_g N_VSS_Mn9@3314_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3315 N_OUT9_Mp9@3315_d N_OUT8_Mp9@3315_g N_VDD_Mp9@3315_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3314 N_OUT9_Mp9@3314_d N_OUT8_Mp9@3314_g N_VDD_Mp9@3314_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3313 N_OUT9_Mn9@3313_d N_OUT8_Mn9@3313_g N_VSS_Mn9@3313_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3312 N_OUT9_Mn9@3312_d N_OUT8_Mn9@3312_g N_VSS_Mn9@3312_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3313 N_OUT9_Mp9@3313_d N_OUT8_Mp9@3313_g N_VDD_Mp9@3313_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3312 N_OUT9_Mp9@3312_d N_OUT8_Mp9@3312_g N_VDD_Mp9@3312_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3311 N_OUT9_Mn9@3311_d N_OUT8_Mn9@3311_g N_VSS_Mn9@3311_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3310 N_OUT9_Mn9@3310_d N_OUT8_Mn9@3310_g N_VSS_Mn9@3310_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3311 N_OUT9_Mp9@3311_d N_OUT8_Mp9@3311_g N_VDD_Mp9@3311_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3310 N_OUT9_Mp9@3310_d N_OUT8_Mp9@3310_g N_VDD_Mp9@3310_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3309 N_OUT9_Mn9@3309_d N_OUT8_Mn9@3309_g N_VSS_Mn9@3309_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3308 N_OUT9_Mn9@3308_d N_OUT8_Mn9@3308_g N_VSS_Mn9@3308_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3309 N_OUT9_Mp9@3309_d N_OUT8_Mp9@3309_g N_VDD_Mp9@3309_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3308 N_OUT9_Mp9@3308_d N_OUT8_Mp9@3308_g N_VDD_Mp9@3308_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3307 N_OUT9_Mn9@3307_d N_OUT8_Mn9@3307_g N_VSS_Mn9@3307_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3306 N_OUT9_Mn9@3306_d N_OUT8_Mn9@3306_g N_VSS_Mn9@3306_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3307 N_OUT9_Mp9@3307_d N_OUT8_Mp9@3307_g N_VDD_Mp9@3307_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3306 N_OUT9_Mp9@3306_d N_OUT8_Mp9@3306_g N_VDD_Mp9@3306_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3305 N_OUT9_Mn9@3305_d N_OUT8_Mn9@3305_g N_VSS_Mn9@3305_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3304 N_OUT9_Mn9@3304_d N_OUT8_Mn9@3304_g N_VSS_Mn9@3304_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3305 N_OUT9_Mp9@3305_d N_OUT8_Mp9@3305_g N_VDD_Mp9@3305_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3304 N_OUT9_Mp9@3304_d N_OUT8_Mp9@3304_g N_VDD_Mp9@3304_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3303 N_OUT9_Mn9@3303_d N_OUT8_Mn9@3303_g N_VSS_Mn9@3303_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3302 N_OUT9_Mn9@3302_d N_OUT8_Mn9@3302_g N_VSS_Mn9@3302_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3303 N_OUT9_Mp9@3303_d N_OUT8_Mp9@3303_g N_VDD_Mp9@3303_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3302 N_OUT9_Mp9@3302_d N_OUT8_Mp9@3302_g N_VDD_Mp9@3302_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3301 N_OUT9_Mn9@3301_d N_OUT8_Mn9@3301_g N_VSS_Mn9@3301_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3300 N_OUT9_Mn9@3300_d N_OUT8_Mn9@3300_g N_VSS_Mn9@3300_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3301 N_OUT9_Mp9@3301_d N_OUT8_Mp9@3301_g N_VDD_Mp9@3301_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3300 N_OUT9_Mp9@3300_d N_OUT8_Mp9@3300_g N_VDD_Mp9@3300_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3299 N_OUT9_Mn9@3299_d N_OUT8_Mn9@3299_g N_VSS_Mn9@3299_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3298 N_OUT9_Mn9@3298_d N_OUT8_Mn9@3298_g N_VSS_Mn9@3298_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3299 N_OUT9_Mp9@3299_d N_OUT8_Mp9@3299_g N_VDD_Mp9@3299_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3298 N_OUT9_Mp9@3298_d N_OUT8_Mp9@3298_g N_VDD_Mp9@3298_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3297 N_OUT9_Mn9@3297_d N_OUT8_Mn9@3297_g N_VSS_Mn9@3297_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3296 N_OUT9_Mn9@3296_d N_OUT8_Mn9@3296_g N_VSS_Mn9@3296_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3297 N_OUT9_Mp9@3297_d N_OUT8_Mp9@3297_g N_VDD_Mp9@3297_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3296 N_OUT9_Mp9@3296_d N_OUT8_Mp9@3296_g N_VDD_Mp9@3296_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3295 N_OUT9_Mn9@3295_d N_OUT8_Mn9@3295_g N_VSS_Mn9@3295_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3294 N_OUT9_Mn9@3294_d N_OUT8_Mn9@3294_g N_VSS_Mn9@3294_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3295 N_OUT9_Mp9@3295_d N_OUT8_Mp9@3295_g N_VDD_Mp9@3295_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3294 N_OUT9_Mp9@3294_d N_OUT8_Mp9@3294_g N_VDD_Mp9@3294_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3293 N_OUT9_Mn9@3293_d N_OUT8_Mn9@3293_g N_VSS_Mn9@3293_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3292 N_OUT9_Mn9@3292_d N_OUT8_Mn9@3292_g N_VSS_Mn9@3292_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3293 N_OUT9_Mp9@3293_d N_OUT8_Mp9@3293_g N_VDD_Mp9@3293_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3292 N_OUT9_Mp9@3292_d N_OUT8_Mp9@3292_g N_VDD_Mp9@3292_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3291 N_OUT9_Mn9@3291_d N_OUT8_Mn9@3291_g N_VSS_Mn9@3291_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3290 N_OUT9_Mn9@3290_d N_OUT8_Mn9@3290_g N_VSS_Mn9@3290_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3291 N_OUT9_Mp9@3291_d N_OUT8_Mp9@3291_g N_VDD_Mp9@3291_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3290 N_OUT9_Mp9@3290_d N_OUT8_Mp9@3290_g N_VDD_Mp9@3290_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3289 N_OUT9_Mn9@3289_d N_OUT8_Mn9@3289_g N_VSS_Mn9@3289_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3288 N_OUT9_Mn9@3288_d N_OUT8_Mn9@3288_g N_VSS_Mn9@3288_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3289 N_OUT9_Mp9@3289_d N_OUT8_Mp9@3289_g N_VDD_Mp9@3289_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3288 N_OUT9_Mp9@3288_d N_OUT8_Mp9@3288_g N_VDD_Mp9@3288_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3287 N_OUT9_Mn9@3287_d N_OUT8_Mn9@3287_g N_VSS_Mn9@3287_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3286 N_OUT9_Mn9@3286_d N_OUT8_Mn9@3286_g N_VSS_Mn9@3286_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3287 N_OUT9_Mp9@3287_d N_OUT8_Mp9@3287_g N_VDD_Mp9@3287_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3286 N_OUT9_Mp9@3286_d N_OUT8_Mp9@3286_g N_VDD_Mp9@3286_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3285 N_OUT9_Mn9@3285_d N_OUT8_Mn9@3285_g N_VSS_Mn9@3285_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3284 N_OUT9_Mn9@3284_d N_OUT8_Mn9@3284_g N_VSS_Mn9@3284_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3285 N_OUT9_Mp9@3285_d N_OUT8_Mp9@3285_g N_VDD_Mp9@3285_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3284 N_OUT9_Mp9@3284_d N_OUT8_Mp9@3284_g N_VDD_Mp9@3284_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3283 N_OUT9_Mn9@3283_d N_OUT8_Mn9@3283_g N_VSS_Mn9@3283_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3282 N_OUT9_Mn9@3282_d N_OUT8_Mn9@3282_g N_VSS_Mn9@3282_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3283 N_OUT9_Mp9@3283_d N_OUT8_Mp9@3283_g N_VDD_Mp9@3283_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3282 N_OUT9_Mp9@3282_d N_OUT8_Mp9@3282_g N_VDD_Mp9@3282_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3281 N_OUT9_Mn9@3281_d N_OUT8_Mn9@3281_g N_VSS_Mn9@3281_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3280 N_OUT9_Mn9@3280_d N_OUT8_Mn9@3280_g N_VSS_Mn9@3280_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3281 N_OUT9_Mp9@3281_d N_OUT8_Mp9@3281_g N_VDD_Mp9@3281_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3280 N_OUT9_Mp9@3280_d N_OUT8_Mp9@3280_g N_VDD_Mp9@3280_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3279 N_OUT9_Mn9@3279_d N_OUT8_Mn9@3279_g N_VSS_Mn9@3279_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3278 N_OUT9_Mn9@3278_d N_OUT8_Mn9@3278_g N_VSS_Mn9@3278_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3279 N_OUT9_Mp9@3279_d N_OUT8_Mp9@3279_g N_VDD_Mp9@3279_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3278 N_OUT9_Mp9@3278_d N_OUT8_Mp9@3278_g N_VDD_Mp9@3278_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3277 N_OUT9_Mn9@3277_d N_OUT8_Mn9@3277_g N_VSS_Mn9@3277_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3276 N_OUT9_Mn9@3276_d N_OUT8_Mn9@3276_g N_VSS_Mn9@3276_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3277 N_OUT9_Mp9@3277_d N_OUT8_Mp9@3277_g N_VDD_Mp9@3277_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3276 N_OUT9_Mp9@3276_d N_OUT8_Mp9@3276_g N_VDD_Mp9@3276_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3275 N_OUT9_Mn9@3275_d N_OUT8_Mn9@3275_g N_VSS_Mn9@3275_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3274 N_OUT9_Mn9@3274_d N_OUT8_Mn9@3274_g N_VSS_Mn9@3274_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3275 N_OUT9_Mp9@3275_d N_OUT8_Mp9@3275_g N_VDD_Mp9@3275_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3274 N_OUT9_Mp9@3274_d N_OUT8_Mp9@3274_g N_VDD_Mp9@3274_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3273 N_OUT9_Mn9@3273_d N_OUT8_Mn9@3273_g N_VSS_Mn9@3273_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3272 N_OUT9_Mn9@3272_d N_OUT8_Mn9@3272_g N_VSS_Mn9@3272_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3273 N_OUT9_Mp9@3273_d N_OUT8_Mp9@3273_g N_VDD_Mp9@3273_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3272 N_OUT9_Mp9@3272_d N_OUT8_Mp9@3272_g N_VDD_Mp9@3272_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3271 N_OUT9_Mn9@3271_d N_OUT8_Mn9@3271_g N_VSS_Mn9@3271_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3270 N_OUT9_Mn9@3270_d N_OUT8_Mn9@3270_g N_VSS_Mn9@3270_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3271 N_OUT9_Mp9@3271_d N_OUT8_Mp9@3271_g N_VDD_Mp9@3271_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3270 N_OUT9_Mp9@3270_d N_OUT8_Mp9@3270_g N_VDD_Mp9@3270_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3269 N_OUT9_Mn9@3269_d N_OUT8_Mn9@3269_g N_VSS_Mn9@3269_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3268 N_OUT9_Mn9@3268_d N_OUT8_Mn9@3268_g N_VSS_Mn9@3268_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3269 N_OUT9_Mp9@3269_d N_OUT8_Mp9@3269_g N_VDD_Mp9@3269_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3268 N_OUT9_Mp9@3268_d N_OUT8_Mp9@3268_g N_VDD_Mp9@3268_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3267 N_OUT9_Mn9@3267_d N_OUT8_Mn9@3267_g N_VSS_Mn9@3267_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3266 N_OUT9_Mn9@3266_d N_OUT8_Mn9@3266_g N_VSS_Mn9@3266_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3267 N_OUT9_Mp9@3267_d N_OUT8_Mp9@3267_g N_VDD_Mp9@3267_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3266 N_OUT9_Mp9@3266_d N_OUT8_Mp9@3266_g N_VDD_Mp9@3266_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3265 N_OUT9_Mn9@3265_d N_OUT8_Mn9@3265_g N_VSS_Mn9@3265_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3264 N_OUT9_Mn9@3264_d N_OUT8_Mn9@3264_g N_VSS_Mn9@3264_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3265 N_OUT9_Mp9@3265_d N_OUT8_Mp9@3265_g N_VDD_Mp9@3265_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3264 N_OUT9_Mp9@3264_d N_OUT8_Mp9@3264_g N_VDD_Mp9@3264_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3263 N_OUT9_Mn9@3263_d N_OUT8_Mn9@3263_g N_VSS_Mn9@3263_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3262 N_OUT9_Mn9@3262_d N_OUT8_Mn9@3262_g N_VSS_Mn9@3262_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3263 N_OUT9_Mp9@3263_d N_OUT8_Mp9@3263_g N_VDD_Mp9@3263_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3262 N_OUT9_Mp9@3262_d N_OUT8_Mp9@3262_g N_VDD_Mp9@3262_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3261 N_OUT9_Mn9@3261_d N_OUT8_Mn9@3261_g N_VSS_Mn9@3261_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3260 N_OUT9_Mn9@3260_d N_OUT8_Mn9@3260_g N_VSS_Mn9@3260_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3261 N_OUT9_Mp9@3261_d N_OUT8_Mp9@3261_g N_VDD_Mp9@3261_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3260 N_OUT9_Mp9@3260_d N_OUT8_Mp9@3260_g N_VDD_Mp9@3260_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3259 N_OUT9_Mn9@3259_d N_OUT8_Mn9@3259_g N_VSS_Mn9@3259_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3258 N_OUT9_Mn9@3258_d N_OUT8_Mn9@3258_g N_VSS_Mn9@3258_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3259 N_OUT9_Mp9@3259_d N_OUT8_Mp9@3259_g N_VDD_Mp9@3259_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3258 N_OUT9_Mp9@3258_d N_OUT8_Mp9@3258_g N_VDD_Mp9@3258_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3257 N_OUT9_Mn9@3257_d N_OUT8_Mn9@3257_g N_VSS_Mn9@3257_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3256 N_OUT9_Mn9@3256_d N_OUT8_Mn9@3256_g N_VSS_Mn9@3256_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3257 N_OUT9_Mp9@3257_d N_OUT8_Mp9@3257_g N_VDD_Mp9@3257_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3256 N_OUT9_Mp9@3256_d N_OUT8_Mp9@3256_g N_VDD_Mp9@3256_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3255 N_OUT9_Mn9@3255_d N_OUT8_Mn9@3255_g N_VSS_Mn9@3255_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3254 N_OUT9_Mn9@3254_d N_OUT8_Mn9@3254_g N_VSS_Mn9@3254_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3255 N_OUT9_Mp9@3255_d N_OUT8_Mp9@3255_g N_VDD_Mp9@3255_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3254 N_OUT9_Mp9@3254_d N_OUT8_Mp9@3254_g N_VDD_Mp9@3254_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3253 N_OUT9_Mn9@3253_d N_OUT8_Mn9@3253_g N_VSS_Mn9@3253_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3252 N_OUT9_Mn9@3252_d N_OUT8_Mn9@3252_g N_VSS_Mn9@3252_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3253 N_OUT9_Mp9@3253_d N_OUT8_Mp9@3253_g N_VDD_Mp9@3253_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3252 N_OUT9_Mp9@3252_d N_OUT8_Mp9@3252_g N_VDD_Mp9@3252_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3251 N_OUT9_Mn9@3251_d N_OUT8_Mn9@3251_g N_VSS_Mn9@3251_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3250 N_OUT9_Mn9@3250_d N_OUT8_Mn9@3250_g N_VSS_Mn9@3250_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3251 N_OUT9_Mp9@3251_d N_OUT8_Mp9@3251_g N_VDD_Mp9@3251_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3250 N_OUT9_Mp9@3250_d N_OUT8_Mp9@3250_g N_VDD_Mp9@3250_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3249 N_OUT9_Mn9@3249_d N_OUT8_Mn9@3249_g N_VSS_Mn9@3249_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3248 N_OUT9_Mn9@3248_d N_OUT8_Mn9@3248_g N_VSS_Mn9@3248_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3249 N_OUT9_Mp9@3249_d N_OUT8_Mp9@3249_g N_VDD_Mp9@3249_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3248 N_OUT9_Mp9@3248_d N_OUT8_Mp9@3248_g N_VDD_Mp9@3248_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3247 N_OUT9_Mn9@3247_d N_OUT8_Mn9@3247_g N_VSS_Mn9@3247_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3246 N_OUT9_Mn9@3246_d N_OUT8_Mn9@3246_g N_VSS_Mn9@3246_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3247 N_OUT9_Mp9@3247_d N_OUT8_Mp9@3247_g N_VDD_Mp9@3247_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3246 N_OUT9_Mp9@3246_d N_OUT8_Mp9@3246_g N_VDD_Mp9@3246_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3245 N_OUT9_Mn9@3245_d N_OUT8_Mn9@3245_g N_VSS_Mn9@3245_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3244 N_OUT9_Mn9@3244_d N_OUT8_Mn9@3244_g N_VSS_Mn9@3244_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3245 N_OUT9_Mp9@3245_d N_OUT8_Mp9@3245_g N_VDD_Mp9@3245_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3244 N_OUT9_Mp9@3244_d N_OUT8_Mp9@3244_g N_VDD_Mp9@3244_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3243 N_OUT9_Mn9@3243_d N_OUT8_Mn9@3243_g N_VSS_Mn9@3243_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3242 N_OUT9_Mn9@3242_d N_OUT8_Mn9@3242_g N_VSS_Mn9@3242_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3243 N_OUT9_Mp9@3243_d N_OUT8_Mp9@3243_g N_VDD_Mp9@3243_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3242 N_OUT9_Mp9@3242_d N_OUT8_Mp9@3242_g N_VDD_Mp9@3242_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3241 N_OUT9_Mn9@3241_d N_OUT8_Mn9@3241_g N_VSS_Mn9@3241_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3240 N_OUT9_Mn9@3240_d N_OUT8_Mn9@3240_g N_VSS_Mn9@3240_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3241 N_OUT9_Mp9@3241_d N_OUT8_Mp9@3241_g N_VDD_Mp9@3241_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3240 N_OUT9_Mp9@3240_d N_OUT8_Mp9@3240_g N_VDD_Mp9@3240_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3239 N_OUT9_Mn9@3239_d N_OUT8_Mn9@3239_g N_VSS_Mn9@3239_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3238 N_OUT9_Mn9@3238_d N_OUT8_Mn9@3238_g N_VSS_Mn9@3238_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3239 N_OUT9_Mp9@3239_d N_OUT8_Mp9@3239_g N_VDD_Mp9@3239_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3238 N_OUT9_Mp9@3238_d N_OUT8_Mp9@3238_g N_VDD_Mp9@3238_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3237 N_OUT9_Mn9@3237_d N_OUT8_Mn9@3237_g N_VSS_Mn9@3237_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3236 N_OUT9_Mn9@3236_d N_OUT8_Mn9@3236_g N_VSS_Mn9@3236_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3237 N_OUT9_Mp9@3237_d N_OUT8_Mp9@3237_g N_VDD_Mp9@3237_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3236 N_OUT9_Mp9@3236_d N_OUT8_Mp9@3236_g N_VDD_Mp9@3236_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3235 N_OUT9_Mn9@3235_d N_OUT8_Mn9@3235_g N_VSS_Mn9@3235_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3234 N_OUT9_Mn9@3234_d N_OUT8_Mn9@3234_g N_VSS_Mn9@3234_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3235 N_OUT9_Mp9@3235_d N_OUT8_Mp9@3235_g N_VDD_Mp9@3235_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3234 N_OUT9_Mp9@3234_d N_OUT8_Mp9@3234_g N_VDD_Mp9@3234_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3233 N_OUT9_Mn9@3233_d N_OUT8_Mn9@3233_g N_VSS_Mn9@3233_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3232 N_OUT9_Mn9@3232_d N_OUT8_Mn9@3232_g N_VSS_Mn9@3232_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3233 N_OUT9_Mp9@3233_d N_OUT8_Mp9@3233_g N_VDD_Mp9@3233_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3232 N_OUT9_Mp9@3232_d N_OUT8_Mp9@3232_g N_VDD_Mp9@3232_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3231 N_OUT9_Mn9@3231_d N_OUT8_Mn9@3231_g N_VSS_Mn9@3231_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3230 N_OUT9_Mn9@3230_d N_OUT8_Mn9@3230_g N_VSS_Mn9@3230_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3231 N_OUT9_Mp9@3231_d N_OUT8_Mp9@3231_g N_VDD_Mp9@3231_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3230 N_OUT9_Mp9@3230_d N_OUT8_Mp9@3230_g N_VDD_Mp9@3230_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3229 N_OUT9_Mn9@3229_d N_OUT8_Mn9@3229_g N_VSS_Mn9@3229_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3228 N_OUT9_Mn9@3228_d N_OUT8_Mn9@3228_g N_VSS_Mn9@3228_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3229 N_OUT9_Mp9@3229_d N_OUT8_Mp9@3229_g N_VDD_Mp9@3229_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3228 N_OUT9_Mp9@3228_d N_OUT8_Mp9@3228_g N_VDD_Mp9@3228_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3227 N_OUT9_Mn9@3227_d N_OUT8_Mn9@3227_g N_VSS_Mn9@3227_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3226 N_OUT9_Mn9@3226_d N_OUT8_Mn9@3226_g N_VSS_Mn9@3226_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3227 N_OUT9_Mp9@3227_d N_OUT8_Mp9@3227_g N_VDD_Mp9@3227_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3226 N_OUT9_Mp9@3226_d N_OUT8_Mp9@3226_g N_VDD_Mp9@3226_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3225 N_OUT9_Mn9@3225_d N_OUT8_Mn9@3225_g N_VSS_Mn9@3225_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3224 N_OUT9_Mn9@3224_d N_OUT8_Mn9@3224_g N_VSS_Mn9@3224_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3225 N_OUT9_Mp9@3225_d N_OUT8_Mp9@3225_g N_VDD_Mp9@3225_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3224 N_OUT9_Mp9@3224_d N_OUT8_Mp9@3224_g N_VDD_Mp9@3224_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3223 N_OUT9_Mn9@3223_d N_OUT8_Mn9@3223_g N_VSS_Mn9@3223_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3222 N_OUT9_Mn9@3222_d N_OUT8_Mn9@3222_g N_VSS_Mn9@3222_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3223 N_OUT9_Mp9@3223_d N_OUT8_Mp9@3223_g N_VDD_Mp9@3223_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3222 N_OUT9_Mp9@3222_d N_OUT8_Mp9@3222_g N_VDD_Mp9@3222_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3221 N_OUT9_Mn9@3221_d N_OUT8_Mn9@3221_g N_VSS_Mn9@3221_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3220 N_OUT9_Mn9@3220_d N_OUT8_Mn9@3220_g N_VSS_Mn9@3220_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3221 N_OUT9_Mp9@3221_d N_OUT8_Mp9@3221_g N_VDD_Mp9@3221_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3220 N_OUT9_Mp9@3220_d N_OUT8_Mp9@3220_g N_VDD_Mp9@3220_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3219 N_OUT9_Mn9@3219_d N_OUT8_Mn9@3219_g N_VSS_Mn9@3219_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3218 N_OUT9_Mn9@3218_d N_OUT8_Mn9@3218_g N_VSS_Mn9@3218_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3219 N_OUT9_Mp9@3219_d N_OUT8_Mp9@3219_g N_VDD_Mp9@3219_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3218 N_OUT9_Mp9@3218_d N_OUT8_Mp9@3218_g N_VDD_Mp9@3218_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3217 N_OUT9_Mn9@3217_d N_OUT8_Mn9@3217_g N_VSS_Mn9@3217_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3216 N_OUT9_Mn9@3216_d N_OUT8_Mn9@3216_g N_VSS_Mn9@3216_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3217 N_OUT9_Mp9@3217_d N_OUT8_Mp9@3217_g N_VDD_Mp9@3217_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3216 N_OUT9_Mp9@3216_d N_OUT8_Mp9@3216_g N_VDD_Mp9@3216_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3215 N_OUT9_Mn9@3215_d N_OUT8_Mn9@3215_g N_VSS_Mn9@3215_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3214 N_OUT9_Mn9@3214_d N_OUT8_Mn9@3214_g N_VSS_Mn9@3214_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3215 N_OUT9_Mp9@3215_d N_OUT8_Mp9@3215_g N_VDD_Mp9@3215_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3214 N_OUT9_Mp9@3214_d N_OUT8_Mp9@3214_g N_VDD_Mp9@3214_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3213 N_OUT9_Mn9@3213_d N_OUT8_Mn9@3213_g N_VSS_Mn9@3213_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3212 N_OUT9_Mn9@3212_d N_OUT8_Mn9@3212_g N_VSS_Mn9@3212_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3213 N_OUT9_Mp9@3213_d N_OUT8_Mp9@3213_g N_VDD_Mp9@3213_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3212 N_OUT9_Mp9@3212_d N_OUT8_Mp9@3212_g N_VDD_Mp9@3212_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3211 N_OUT9_Mn9@3211_d N_OUT8_Mn9@3211_g N_VSS_Mn9@3211_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3210 N_OUT9_Mn9@3210_d N_OUT8_Mn9@3210_g N_VSS_Mn9@3210_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3211 N_OUT9_Mp9@3211_d N_OUT8_Mp9@3211_g N_VDD_Mp9@3211_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3210 N_OUT9_Mp9@3210_d N_OUT8_Mp9@3210_g N_VDD_Mp9@3210_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3209 N_OUT9_Mn9@3209_d N_OUT8_Mn9@3209_g N_VSS_Mn9@3209_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3208 N_OUT9_Mn9@3208_d N_OUT8_Mn9@3208_g N_VSS_Mn9@3208_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3209 N_OUT9_Mp9@3209_d N_OUT8_Mp9@3209_g N_VDD_Mp9@3209_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3208 N_OUT9_Mp9@3208_d N_OUT8_Mp9@3208_g N_VDD_Mp9@3208_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3207 N_OUT9_Mn9@3207_d N_OUT8_Mn9@3207_g N_VSS_Mn9@3207_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3206 N_OUT9_Mn9@3206_d N_OUT8_Mn9@3206_g N_VSS_Mn9@3206_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3207 N_OUT9_Mp9@3207_d N_OUT8_Mp9@3207_g N_VDD_Mp9@3207_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3206 N_OUT9_Mp9@3206_d N_OUT8_Mp9@3206_g N_VDD_Mp9@3206_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3205 N_OUT9_Mn9@3205_d N_OUT8_Mn9@3205_g N_VSS_Mn9@3205_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3204 N_OUT9_Mn9@3204_d N_OUT8_Mn9@3204_g N_VSS_Mn9@3204_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3205 N_OUT9_Mp9@3205_d N_OUT8_Mp9@3205_g N_VDD_Mp9@3205_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3204 N_OUT9_Mp9@3204_d N_OUT8_Mp9@3204_g N_VDD_Mp9@3204_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3203 N_OUT9_Mn9@3203_d N_OUT8_Mn9@3203_g N_VSS_Mn9@3203_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3202 N_OUT9_Mn9@3202_d N_OUT8_Mn9@3202_g N_VSS_Mn9@3202_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3203 N_OUT9_Mp9@3203_d N_OUT8_Mp9@3203_g N_VDD_Mp9@3203_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3202 N_OUT9_Mp9@3202_d N_OUT8_Mp9@3202_g N_VDD_Mp9@3202_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3201 N_OUT9_Mn9@3201_d N_OUT8_Mn9@3201_g N_VSS_Mn9@3201_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3200 N_OUT9_Mn9@3200_d N_OUT8_Mn9@3200_g N_VSS_Mn9@3200_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3201 N_OUT9_Mp9@3201_d N_OUT8_Mp9@3201_g N_VDD_Mp9@3201_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3200 N_OUT9_Mp9@3200_d N_OUT8_Mp9@3200_g N_VDD_Mp9@3200_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3199 N_OUT9_Mn9@3199_d N_OUT8_Mn9@3199_g N_VSS_Mn9@3199_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3198 N_OUT9_Mn9@3198_d N_OUT8_Mn9@3198_g N_VSS_Mn9@3198_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3199 N_OUT9_Mp9@3199_d N_OUT8_Mp9@3199_g N_VDD_Mp9@3199_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3198 N_OUT9_Mp9@3198_d N_OUT8_Mp9@3198_g N_VDD_Mp9@3198_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3197 N_OUT9_Mn9@3197_d N_OUT8_Mn9@3197_g N_VSS_Mn9@3197_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3196 N_OUT9_Mn9@3196_d N_OUT8_Mn9@3196_g N_VSS_Mn9@3196_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3197 N_OUT9_Mp9@3197_d N_OUT8_Mp9@3197_g N_VDD_Mp9@3197_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3196 N_OUT9_Mp9@3196_d N_OUT8_Mp9@3196_g N_VDD_Mp9@3196_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3195 N_OUT9_Mn9@3195_d N_OUT8_Mn9@3195_g N_VSS_Mn9@3195_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3194 N_OUT9_Mn9@3194_d N_OUT8_Mn9@3194_g N_VSS_Mn9@3194_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3195 N_OUT9_Mp9@3195_d N_OUT8_Mp9@3195_g N_VDD_Mp9@3195_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3194 N_OUT9_Mp9@3194_d N_OUT8_Mp9@3194_g N_VDD_Mp9@3194_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3193 N_OUT9_Mn9@3193_d N_OUT8_Mn9@3193_g N_VSS_Mn9@3193_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3192 N_OUT9_Mn9@3192_d N_OUT8_Mn9@3192_g N_VSS_Mn9@3192_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3193 N_OUT9_Mp9@3193_d N_OUT8_Mp9@3193_g N_VDD_Mp9@3193_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3192 N_OUT9_Mp9@3192_d N_OUT8_Mp9@3192_g N_VDD_Mp9@3192_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3191 N_OUT9_Mn9@3191_d N_OUT8_Mn9@3191_g N_VSS_Mn9@3191_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3190 N_OUT9_Mn9@3190_d N_OUT8_Mn9@3190_g N_VSS_Mn9@3190_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3191 N_OUT9_Mp9@3191_d N_OUT8_Mp9@3191_g N_VDD_Mp9@3191_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3190 N_OUT9_Mp9@3190_d N_OUT8_Mp9@3190_g N_VDD_Mp9@3190_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3189 N_OUT9_Mn9@3189_d N_OUT8_Mn9@3189_g N_VSS_Mn9@3189_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3188 N_OUT9_Mn9@3188_d N_OUT8_Mn9@3188_g N_VSS_Mn9@3188_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3189 N_OUT9_Mp9@3189_d N_OUT8_Mp9@3189_g N_VDD_Mp9@3189_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3188 N_OUT9_Mp9@3188_d N_OUT8_Mp9@3188_g N_VDD_Mp9@3188_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3187 N_OUT9_Mn9@3187_d N_OUT8_Mn9@3187_g N_VSS_Mn9@3187_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3186 N_OUT9_Mn9@3186_d N_OUT8_Mn9@3186_g N_VSS_Mn9@3186_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3187 N_OUT9_Mp9@3187_d N_OUT8_Mp9@3187_g N_VDD_Mp9@3187_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3186 N_OUT9_Mp9@3186_d N_OUT8_Mp9@3186_g N_VDD_Mp9@3186_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3185 N_OUT9_Mn9@3185_d N_OUT8_Mn9@3185_g N_VSS_Mn9@3185_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3184 N_OUT9_Mn9@3184_d N_OUT8_Mn9@3184_g N_VSS_Mn9@3184_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3185 N_OUT9_Mp9@3185_d N_OUT8_Mp9@3185_g N_VDD_Mp9@3185_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3184 N_OUT9_Mp9@3184_d N_OUT8_Mp9@3184_g N_VDD_Mp9@3184_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3183 N_OUT9_Mn9@3183_d N_OUT8_Mn9@3183_g N_VSS_Mn9@3183_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3182 N_OUT9_Mn9@3182_d N_OUT8_Mn9@3182_g N_VSS_Mn9@3182_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3183 N_OUT9_Mp9@3183_d N_OUT8_Mp9@3183_g N_VDD_Mp9@3183_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3182 N_OUT9_Mp9@3182_d N_OUT8_Mp9@3182_g N_VDD_Mp9@3182_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3181 N_OUT9_Mn9@3181_d N_OUT8_Mn9@3181_g N_VSS_Mn9@3181_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3180 N_OUT9_Mn9@3180_d N_OUT8_Mn9@3180_g N_VSS_Mn9@3180_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3181 N_OUT9_Mp9@3181_d N_OUT8_Mp9@3181_g N_VDD_Mp9@3181_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3180 N_OUT9_Mp9@3180_d N_OUT8_Mp9@3180_g N_VDD_Mp9@3180_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3179 N_OUT9_Mn9@3179_d N_OUT8_Mn9@3179_g N_VSS_Mn9@3179_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3178 N_OUT9_Mn9@3178_d N_OUT8_Mn9@3178_g N_VSS_Mn9@3178_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3179 N_OUT9_Mp9@3179_d N_OUT8_Mp9@3179_g N_VDD_Mp9@3179_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3178 N_OUT9_Mp9@3178_d N_OUT8_Mp9@3178_g N_VDD_Mp9@3178_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3177 N_OUT9_Mn9@3177_d N_OUT8_Mn9@3177_g N_VSS_Mn9@3177_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3176 N_OUT9_Mn9@3176_d N_OUT8_Mn9@3176_g N_VSS_Mn9@3176_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3177 N_OUT9_Mp9@3177_d N_OUT8_Mp9@3177_g N_VDD_Mp9@3177_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3176 N_OUT9_Mp9@3176_d N_OUT8_Mp9@3176_g N_VDD_Mp9@3176_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3175 N_OUT9_Mn9@3175_d N_OUT8_Mn9@3175_g N_VSS_Mn9@3175_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3174 N_OUT9_Mn9@3174_d N_OUT8_Mn9@3174_g N_VSS_Mn9@3174_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3175 N_OUT9_Mp9@3175_d N_OUT8_Mp9@3175_g N_VDD_Mp9@3175_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3174 N_OUT9_Mp9@3174_d N_OUT8_Mp9@3174_g N_VDD_Mp9@3174_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3173 N_OUT9_Mn9@3173_d N_OUT8_Mn9@3173_g N_VSS_Mn9@3173_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3172 N_OUT9_Mn9@3172_d N_OUT8_Mn9@3172_g N_VSS_Mn9@3172_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3173 N_OUT9_Mp9@3173_d N_OUT8_Mp9@3173_g N_VDD_Mp9@3173_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3172 N_OUT9_Mp9@3172_d N_OUT8_Mp9@3172_g N_VDD_Mp9@3172_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3171 N_OUT9_Mn9@3171_d N_OUT8_Mn9@3171_g N_VSS_Mn9@3171_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3170 N_OUT9_Mn9@3170_d N_OUT8_Mn9@3170_g N_VSS_Mn9@3170_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3171 N_OUT9_Mp9@3171_d N_OUT8_Mp9@3171_g N_VDD_Mp9@3171_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3170 N_OUT9_Mp9@3170_d N_OUT8_Mp9@3170_g N_VDD_Mp9@3170_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3169 N_OUT9_Mn9@3169_d N_OUT8_Mn9@3169_g N_VSS_Mn9@3169_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3168 N_OUT9_Mn9@3168_d N_OUT8_Mn9@3168_g N_VSS_Mn9@3168_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3169 N_OUT9_Mp9@3169_d N_OUT8_Mp9@3169_g N_VDD_Mp9@3169_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3168 N_OUT9_Mp9@3168_d N_OUT8_Mp9@3168_g N_VDD_Mp9@3168_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3167 N_OUT9_Mn9@3167_d N_OUT8_Mn9@3167_g N_VSS_Mn9@3167_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3166 N_OUT9_Mn9@3166_d N_OUT8_Mn9@3166_g N_VSS_Mn9@3166_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3167 N_OUT9_Mp9@3167_d N_OUT8_Mp9@3167_g N_VDD_Mp9@3167_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3166 N_OUT9_Mp9@3166_d N_OUT8_Mp9@3166_g N_VDD_Mp9@3166_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3165 N_OUT9_Mn9@3165_d N_OUT8_Mn9@3165_g N_VSS_Mn9@3165_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3164 N_OUT9_Mn9@3164_d N_OUT8_Mn9@3164_g N_VSS_Mn9@3164_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3165 N_OUT9_Mp9@3165_d N_OUT8_Mp9@3165_g N_VDD_Mp9@3165_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3164 N_OUT9_Mp9@3164_d N_OUT8_Mp9@3164_g N_VDD_Mp9@3164_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3163 N_OUT9_Mn9@3163_d N_OUT8_Mn9@3163_g N_VSS_Mn9@3163_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3162 N_OUT9_Mn9@3162_d N_OUT8_Mn9@3162_g N_VSS_Mn9@3162_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3163 N_OUT9_Mp9@3163_d N_OUT8_Mp9@3163_g N_VDD_Mp9@3163_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3162 N_OUT9_Mp9@3162_d N_OUT8_Mp9@3162_g N_VDD_Mp9@3162_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3161 N_OUT9_Mn9@3161_d N_OUT8_Mn9@3161_g N_VSS_Mn9@3161_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3160 N_OUT9_Mn9@3160_d N_OUT8_Mn9@3160_g N_VSS_Mn9@3160_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3161 N_OUT9_Mp9@3161_d N_OUT8_Mp9@3161_g N_VDD_Mp9@3161_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3160 N_OUT9_Mp9@3160_d N_OUT8_Mp9@3160_g N_VDD_Mp9@3160_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3159 N_OUT9_Mn9@3159_d N_OUT8_Mn9@3159_g N_VSS_Mn9@3159_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3158 N_OUT9_Mn9@3158_d N_OUT8_Mn9@3158_g N_VSS_Mn9@3158_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3159 N_OUT9_Mp9@3159_d N_OUT8_Mp9@3159_g N_VDD_Mp9@3159_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3158 N_OUT9_Mp9@3158_d N_OUT8_Mp9@3158_g N_VDD_Mp9@3158_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3157 N_OUT9_Mn9@3157_d N_OUT8_Mn9@3157_g N_VSS_Mn9@3157_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3156 N_OUT9_Mn9@3156_d N_OUT8_Mn9@3156_g N_VSS_Mn9@3156_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3157 N_OUT9_Mp9@3157_d N_OUT8_Mp9@3157_g N_VDD_Mp9@3157_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3156 N_OUT9_Mp9@3156_d N_OUT8_Mp9@3156_g N_VDD_Mp9@3156_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3155 N_OUT9_Mn9@3155_d N_OUT8_Mn9@3155_g N_VSS_Mn9@3155_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3154 N_OUT9_Mn9@3154_d N_OUT8_Mn9@3154_g N_VSS_Mn9@3154_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3155 N_OUT9_Mp9@3155_d N_OUT8_Mp9@3155_g N_VDD_Mp9@3155_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3154 N_OUT9_Mp9@3154_d N_OUT8_Mp9@3154_g N_VDD_Mp9@3154_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3153 N_OUT9_Mn9@3153_d N_OUT8_Mn9@3153_g N_VSS_Mn9@3153_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3152 N_OUT9_Mn9@3152_d N_OUT8_Mn9@3152_g N_VSS_Mn9@3152_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3153 N_OUT9_Mp9@3153_d N_OUT8_Mp9@3153_g N_VDD_Mp9@3153_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3152 N_OUT9_Mp9@3152_d N_OUT8_Mp9@3152_g N_VDD_Mp9@3152_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3151 N_OUT9_Mn9@3151_d N_OUT8_Mn9@3151_g N_VSS_Mn9@3151_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3150 N_OUT9_Mn9@3150_d N_OUT8_Mn9@3150_g N_VSS_Mn9@3150_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3151 N_OUT9_Mp9@3151_d N_OUT8_Mp9@3151_g N_VDD_Mp9@3151_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3150 N_OUT9_Mp9@3150_d N_OUT8_Mp9@3150_g N_VDD_Mp9@3150_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3149 N_OUT9_Mn9@3149_d N_OUT8_Mn9@3149_g N_VSS_Mn9@3149_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3148 N_OUT9_Mn9@3148_d N_OUT8_Mn9@3148_g N_VSS_Mn9@3148_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3149 N_OUT9_Mp9@3149_d N_OUT8_Mp9@3149_g N_VDD_Mp9@3149_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3148 N_OUT9_Mp9@3148_d N_OUT8_Mp9@3148_g N_VDD_Mp9@3148_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3147 N_OUT9_Mn9@3147_d N_OUT8_Mn9@3147_g N_VSS_Mn9@3147_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3146 N_OUT9_Mn9@3146_d N_OUT8_Mn9@3146_g N_VSS_Mn9@3146_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3147 N_OUT9_Mp9@3147_d N_OUT8_Mp9@3147_g N_VDD_Mp9@3147_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3146 N_OUT9_Mp9@3146_d N_OUT8_Mp9@3146_g N_VDD_Mp9@3146_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3145 N_OUT9_Mn9@3145_d N_OUT8_Mn9@3145_g N_VSS_Mn9@3145_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3144 N_OUT9_Mn9@3144_d N_OUT8_Mn9@3144_g N_VSS_Mn9@3144_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3145 N_OUT9_Mp9@3145_d N_OUT8_Mp9@3145_g N_VDD_Mp9@3145_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3144 N_OUT9_Mp9@3144_d N_OUT8_Mp9@3144_g N_VDD_Mp9@3144_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3143 N_OUT9_Mn9@3143_d N_OUT8_Mn9@3143_g N_VSS_Mn9@3143_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3142 N_OUT9_Mn9@3142_d N_OUT8_Mn9@3142_g N_VSS_Mn9@3142_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3143 N_OUT9_Mp9@3143_d N_OUT8_Mp9@3143_g N_VDD_Mp9@3143_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3142 N_OUT9_Mp9@3142_d N_OUT8_Mp9@3142_g N_VDD_Mp9@3142_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3141 N_OUT9_Mn9@3141_d N_OUT8_Mn9@3141_g N_VSS_Mn9@3141_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3140 N_OUT9_Mn9@3140_d N_OUT8_Mn9@3140_g N_VSS_Mn9@3140_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3141 N_OUT9_Mp9@3141_d N_OUT8_Mp9@3141_g N_VDD_Mp9@3141_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3140 N_OUT9_Mp9@3140_d N_OUT8_Mp9@3140_g N_VDD_Mp9@3140_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3139 N_OUT9_Mn9@3139_d N_OUT8_Mn9@3139_g N_VSS_Mn9@3139_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3138 N_OUT9_Mn9@3138_d N_OUT8_Mn9@3138_g N_VSS_Mn9@3138_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3139 N_OUT9_Mp9@3139_d N_OUT8_Mp9@3139_g N_VDD_Mp9@3139_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3138 N_OUT9_Mp9@3138_d N_OUT8_Mp9@3138_g N_VDD_Mp9@3138_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3137 N_OUT9_Mn9@3137_d N_OUT8_Mn9@3137_g N_VSS_Mn9@3137_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3136 N_OUT9_Mn9@3136_d N_OUT8_Mn9@3136_g N_VSS_Mn9@3136_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3137 N_OUT9_Mp9@3137_d N_OUT8_Mp9@3137_g N_VDD_Mp9@3137_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3136 N_OUT9_Mp9@3136_d N_OUT8_Mp9@3136_g N_VDD_Mp9@3136_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3135 N_OUT9_Mn9@3135_d N_OUT8_Mn9@3135_g N_VSS_Mn9@3135_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3134 N_OUT9_Mn9@3134_d N_OUT8_Mn9@3134_g N_VSS_Mn9@3134_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3135 N_OUT9_Mp9@3135_d N_OUT8_Mp9@3135_g N_VDD_Mp9@3135_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3134 N_OUT9_Mp9@3134_d N_OUT8_Mp9@3134_g N_VDD_Mp9@3134_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3133 N_OUT9_Mn9@3133_d N_OUT8_Mn9@3133_g N_VSS_Mn9@3133_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3132 N_OUT9_Mn9@3132_d N_OUT8_Mn9@3132_g N_VSS_Mn9@3132_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3133 N_OUT9_Mp9@3133_d N_OUT8_Mp9@3133_g N_VDD_Mp9@3133_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3132 N_OUT9_Mp9@3132_d N_OUT8_Mp9@3132_g N_VDD_Mp9@3132_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3131 N_OUT9_Mn9@3131_d N_OUT8_Mn9@3131_g N_VSS_Mn9@3131_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3130 N_OUT9_Mn9@3130_d N_OUT8_Mn9@3130_g N_VSS_Mn9@3130_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3131 N_OUT9_Mp9@3131_d N_OUT8_Mp9@3131_g N_VDD_Mp9@3131_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3130 N_OUT9_Mp9@3130_d N_OUT8_Mp9@3130_g N_VDD_Mp9@3130_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3129 N_OUT9_Mn9@3129_d N_OUT8_Mn9@3129_g N_VSS_Mn9@3129_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3128 N_OUT9_Mn9@3128_d N_OUT8_Mn9@3128_g N_VSS_Mn9@3128_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3129 N_OUT9_Mp9@3129_d N_OUT8_Mp9@3129_g N_VDD_Mp9@3129_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3128 N_OUT9_Mp9@3128_d N_OUT8_Mp9@3128_g N_VDD_Mp9@3128_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3127 N_OUT9_Mn9@3127_d N_OUT8_Mn9@3127_g N_VSS_Mn9@3127_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3126 N_OUT9_Mn9@3126_d N_OUT8_Mn9@3126_g N_VSS_Mn9@3126_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3127 N_OUT9_Mp9@3127_d N_OUT8_Mp9@3127_g N_VDD_Mp9@3127_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3126 N_OUT9_Mp9@3126_d N_OUT8_Mp9@3126_g N_VDD_Mp9@3126_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3125 N_OUT9_Mn9@3125_d N_OUT8_Mn9@3125_g N_VSS_Mn9@3125_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3124 N_OUT9_Mn9@3124_d N_OUT8_Mn9@3124_g N_VSS_Mn9@3124_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3125 N_OUT9_Mp9@3125_d N_OUT8_Mp9@3125_g N_VDD_Mp9@3125_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3124 N_OUT9_Mp9@3124_d N_OUT8_Mp9@3124_g N_VDD_Mp9@3124_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3123 N_OUT9_Mn9@3123_d N_OUT8_Mn9@3123_g N_VSS_Mn9@3123_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3122 N_OUT9_Mn9@3122_d N_OUT8_Mn9@3122_g N_VSS_Mn9@3122_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3123 N_OUT9_Mp9@3123_d N_OUT8_Mp9@3123_g N_VDD_Mp9@3123_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3122 N_OUT9_Mp9@3122_d N_OUT8_Mp9@3122_g N_VDD_Mp9@3122_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3121 N_OUT9_Mn9@3121_d N_OUT8_Mn9@3121_g N_VSS_Mn9@3121_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3120 N_OUT9_Mn9@3120_d N_OUT8_Mn9@3120_g N_VSS_Mn9@3120_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3121 N_OUT9_Mp9@3121_d N_OUT8_Mp9@3121_g N_VDD_Mp9@3121_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3120 N_OUT9_Mp9@3120_d N_OUT8_Mp9@3120_g N_VDD_Mp9@3120_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3119 N_OUT9_Mn9@3119_d N_OUT8_Mn9@3119_g N_VSS_Mn9@3119_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3118 N_OUT9_Mn9@3118_d N_OUT8_Mn9@3118_g N_VSS_Mn9@3118_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3119 N_OUT9_Mp9@3119_d N_OUT8_Mp9@3119_g N_VDD_Mp9@3119_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3118 N_OUT9_Mp9@3118_d N_OUT8_Mp9@3118_g N_VDD_Mp9@3118_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3117 N_OUT9_Mn9@3117_d N_OUT8_Mn9@3117_g N_VSS_Mn9@3117_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3116 N_OUT9_Mn9@3116_d N_OUT8_Mn9@3116_g N_VSS_Mn9@3116_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3117 N_OUT9_Mp9@3117_d N_OUT8_Mp9@3117_g N_VDD_Mp9@3117_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3116 N_OUT9_Mp9@3116_d N_OUT8_Mp9@3116_g N_VDD_Mp9@3116_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3115 N_OUT9_Mn9@3115_d N_OUT8_Mn9@3115_g N_VSS_Mn9@3115_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3114 N_OUT9_Mn9@3114_d N_OUT8_Mn9@3114_g N_VSS_Mn9@3114_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3115 N_OUT9_Mp9@3115_d N_OUT8_Mp9@3115_g N_VDD_Mp9@3115_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3114 N_OUT9_Mp9@3114_d N_OUT8_Mp9@3114_g N_VDD_Mp9@3114_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3113 N_OUT9_Mn9@3113_d N_OUT8_Mn9@3113_g N_VSS_Mn9@3113_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3112 N_OUT9_Mn9@3112_d N_OUT8_Mn9@3112_g N_VSS_Mn9@3112_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3113 N_OUT9_Mp9@3113_d N_OUT8_Mp9@3113_g N_VDD_Mp9@3113_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3112 N_OUT9_Mp9@3112_d N_OUT8_Mp9@3112_g N_VDD_Mp9@3112_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3111 N_OUT9_Mn9@3111_d N_OUT8_Mn9@3111_g N_VSS_Mn9@3111_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3110 N_OUT9_Mn9@3110_d N_OUT8_Mn9@3110_g N_VSS_Mn9@3110_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3111 N_OUT9_Mp9@3111_d N_OUT8_Mp9@3111_g N_VDD_Mp9@3111_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3110 N_OUT9_Mp9@3110_d N_OUT8_Mp9@3110_g N_VDD_Mp9@3110_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3109 N_OUT9_Mn9@3109_d N_OUT8_Mn9@3109_g N_VSS_Mn9@3109_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3108 N_OUT9_Mn9@3108_d N_OUT8_Mn9@3108_g N_VSS_Mn9@3108_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3109 N_OUT9_Mp9@3109_d N_OUT8_Mp9@3109_g N_VDD_Mp9@3109_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3108 N_OUT9_Mp9@3108_d N_OUT8_Mp9@3108_g N_VDD_Mp9@3108_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3107 N_OUT9_Mn9@3107_d N_OUT8_Mn9@3107_g N_VSS_Mn9@3107_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3106 N_OUT9_Mn9@3106_d N_OUT8_Mn9@3106_g N_VSS_Mn9@3106_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3107 N_OUT9_Mp9@3107_d N_OUT8_Mp9@3107_g N_VDD_Mp9@3107_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3106 N_OUT9_Mp9@3106_d N_OUT8_Mp9@3106_g N_VDD_Mp9@3106_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3105 N_OUT9_Mn9@3105_d N_OUT8_Mn9@3105_g N_VSS_Mn9@3105_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3104 N_OUT9_Mn9@3104_d N_OUT8_Mn9@3104_g N_VSS_Mn9@3104_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3105 N_OUT9_Mp9@3105_d N_OUT8_Mp9@3105_g N_VDD_Mp9@3105_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3104 N_OUT9_Mp9@3104_d N_OUT8_Mp9@3104_g N_VDD_Mp9@3104_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3103 N_OUT9_Mn9@3103_d N_OUT8_Mn9@3103_g N_VSS_Mn9@3103_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3102 N_OUT9_Mn9@3102_d N_OUT8_Mn9@3102_g N_VSS_Mn9@3102_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3103 N_OUT9_Mp9@3103_d N_OUT8_Mp9@3103_g N_VDD_Mp9@3103_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3102 N_OUT9_Mp9@3102_d N_OUT8_Mp9@3102_g N_VDD_Mp9@3102_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3101 N_OUT9_Mn9@3101_d N_OUT8_Mn9@3101_g N_VSS_Mn9@3101_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3100 N_OUT9_Mn9@3100_d N_OUT8_Mn9@3100_g N_VSS_Mn9@3100_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3101 N_OUT9_Mp9@3101_d N_OUT8_Mp9@3101_g N_VDD_Mp9@3101_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3100 N_OUT9_Mp9@3100_d N_OUT8_Mp9@3100_g N_VDD_Mp9@3100_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3099 N_OUT9_Mn9@3099_d N_OUT8_Mn9@3099_g N_VSS_Mn9@3099_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3098 N_OUT9_Mn9@3098_d N_OUT8_Mn9@3098_g N_VSS_Mn9@3098_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3099 N_OUT9_Mp9@3099_d N_OUT8_Mp9@3099_g N_VDD_Mp9@3099_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3098 N_OUT9_Mp9@3098_d N_OUT8_Mp9@3098_g N_VDD_Mp9@3098_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3097 N_OUT9_Mn9@3097_d N_OUT8_Mn9@3097_g N_VSS_Mn9@3097_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3096 N_OUT9_Mn9@3096_d N_OUT8_Mn9@3096_g N_VSS_Mn9@3096_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3097 N_OUT9_Mp9@3097_d N_OUT8_Mp9@3097_g N_VDD_Mp9@3097_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3096 N_OUT9_Mp9@3096_d N_OUT8_Mp9@3096_g N_VDD_Mp9@3096_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3095 N_OUT9_Mn9@3095_d N_OUT8_Mn9@3095_g N_VSS_Mn9@3095_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3094 N_OUT9_Mn9@3094_d N_OUT8_Mn9@3094_g N_VSS_Mn9@3094_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3095 N_OUT9_Mp9@3095_d N_OUT8_Mp9@3095_g N_VDD_Mp9@3095_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3094 N_OUT9_Mp9@3094_d N_OUT8_Mp9@3094_g N_VDD_Mp9@3094_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3093 N_OUT9_Mn9@3093_d N_OUT8_Mn9@3093_g N_VSS_Mn9@3093_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3092 N_OUT9_Mn9@3092_d N_OUT8_Mn9@3092_g N_VSS_Mn9@3092_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3093 N_OUT9_Mp9@3093_d N_OUT8_Mp9@3093_g N_VDD_Mp9@3093_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3092 N_OUT9_Mp9@3092_d N_OUT8_Mp9@3092_g N_VDD_Mp9@3092_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3091 N_OUT9_Mn9@3091_d N_OUT8_Mn9@3091_g N_VSS_Mn9@3091_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3090 N_OUT9_Mn9@3090_d N_OUT8_Mn9@3090_g N_VSS_Mn9@3090_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3091 N_OUT9_Mp9@3091_d N_OUT8_Mp9@3091_g N_VDD_Mp9@3091_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3090 N_OUT9_Mp9@3090_d N_OUT8_Mp9@3090_g N_VDD_Mp9@3090_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3089 N_OUT9_Mn9@3089_d N_OUT8_Mn9@3089_g N_VSS_Mn9@3089_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3088 N_OUT9_Mn9@3088_d N_OUT8_Mn9@3088_g N_VSS_Mn9@3088_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3089 N_OUT9_Mp9@3089_d N_OUT8_Mp9@3089_g N_VDD_Mp9@3089_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3088 N_OUT9_Mp9@3088_d N_OUT8_Mp9@3088_g N_VDD_Mp9@3088_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3087 N_OUT9_Mn9@3087_d N_OUT8_Mn9@3087_g N_VSS_Mn9@3087_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3086 N_OUT9_Mn9@3086_d N_OUT8_Mn9@3086_g N_VSS_Mn9@3086_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3087 N_OUT9_Mp9@3087_d N_OUT8_Mp9@3087_g N_VDD_Mp9@3087_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3086 N_OUT9_Mp9@3086_d N_OUT8_Mp9@3086_g N_VDD_Mp9@3086_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3085 N_OUT9_Mn9@3085_d N_OUT8_Mn9@3085_g N_VSS_Mn9@3085_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3084 N_OUT9_Mn9@3084_d N_OUT8_Mn9@3084_g N_VSS_Mn9@3084_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3085 N_OUT9_Mp9@3085_d N_OUT8_Mp9@3085_g N_VDD_Mp9@3085_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3084 N_OUT9_Mp9@3084_d N_OUT8_Mp9@3084_g N_VDD_Mp9@3084_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3083 N_OUT9_Mn9@3083_d N_OUT8_Mn9@3083_g N_VSS_Mn9@3083_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3082 N_OUT9_Mn9@3082_d N_OUT8_Mn9@3082_g N_VSS_Mn9@3082_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3083 N_OUT9_Mp9@3083_d N_OUT8_Mp9@3083_g N_VDD_Mp9@3083_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3082 N_OUT9_Mp9@3082_d N_OUT8_Mp9@3082_g N_VDD_Mp9@3082_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3081 N_OUT9_Mn9@3081_d N_OUT8_Mn9@3081_g N_VSS_Mn9@3081_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3080 N_OUT9_Mn9@3080_d N_OUT8_Mn9@3080_g N_VSS_Mn9@3080_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3081 N_OUT9_Mp9@3081_d N_OUT8_Mp9@3081_g N_VDD_Mp9@3081_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3080 N_OUT9_Mp9@3080_d N_OUT8_Mp9@3080_g N_VDD_Mp9@3080_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3079 N_OUT9_Mn9@3079_d N_OUT8_Mn9@3079_g N_VSS_Mn9@3079_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3078 N_OUT9_Mn9@3078_d N_OUT8_Mn9@3078_g N_VSS_Mn9@3078_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3079 N_OUT9_Mp9@3079_d N_OUT8_Mp9@3079_g N_VDD_Mp9@3079_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3078 N_OUT9_Mp9@3078_d N_OUT8_Mp9@3078_g N_VDD_Mp9@3078_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3077 N_OUT9_Mn9@3077_d N_OUT8_Mn9@3077_g N_VSS_Mn9@3077_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3076 N_OUT9_Mn9@3076_d N_OUT8_Mn9@3076_g N_VSS_Mn9@3076_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3077 N_OUT9_Mp9@3077_d N_OUT8_Mp9@3077_g N_VDD_Mp9@3077_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3076 N_OUT9_Mp9@3076_d N_OUT8_Mp9@3076_g N_VDD_Mp9@3076_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3075 N_OUT9_Mn9@3075_d N_OUT8_Mn9@3075_g N_VSS_Mn9@3075_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3074 N_OUT9_Mn9@3074_d N_OUT8_Mn9@3074_g N_VSS_Mn9@3074_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3075 N_OUT9_Mp9@3075_d N_OUT8_Mp9@3075_g N_VDD_Mp9@3075_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3074 N_OUT9_Mp9@3074_d N_OUT8_Mp9@3074_g N_VDD_Mp9@3074_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3073 N_OUT9_Mn9@3073_d N_OUT8_Mn9@3073_g N_VSS_Mn9@3073_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3072 N_OUT9_Mn9@3072_d N_OUT8_Mn9@3072_g N_VSS_Mn9@3072_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3073 N_OUT9_Mp9@3073_d N_OUT8_Mp9@3073_g N_VDD_Mp9@3073_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3072 N_OUT9_Mp9@3072_d N_OUT8_Mp9@3072_g N_VDD_Mp9@3072_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3071 N_OUT9_Mn9@3071_d N_OUT8_Mn9@3071_g N_VSS_Mn9@3071_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3070 N_OUT9_Mn9@3070_d N_OUT8_Mn9@3070_g N_VSS_Mn9@3070_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3071 N_OUT9_Mp9@3071_d N_OUT8_Mp9@3071_g N_VDD_Mp9@3071_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3070 N_OUT9_Mp9@3070_d N_OUT8_Mp9@3070_g N_VDD_Mp9@3070_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3069 N_OUT9_Mn9@3069_d N_OUT8_Mn9@3069_g N_VSS_Mn9@3069_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3068 N_OUT9_Mn9@3068_d N_OUT8_Mn9@3068_g N_VSS_Mn9@3068_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3069 N_OUT9_Mp9@3069_d N_OUT8_Mp9@3069_g N_VDD_Mp9@3069_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3068 N_OUT9_Mp9@3068_d N_OUT8_Mp9@3068_g N_VDD_Mp9@3068_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3067 N_OUT9_Mn9@3067_d N_OUT8_Mn9@3067_g N_VSS_Mn9@3067_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3066 N_OUT9_Mn9@3066_d N_OUT8_Mn9@3066_g N_VSS_Mn9@3066_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3067 N_OUT9_Mp9@3067_d N_OUT8_Mp9@3067_g N_VDD_Mp9@3067_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3066 N_OUT9_Mp9@3066_d N_OUT8_Mp9@3066_g N_VDD_Mp9@3066_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3065 N_OUT9_Mn9@3065_d N_OUT8_Mn9@3065_g N_VSS_Mn9@3065_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3064 N_OUT9_Mn9@3064_d N_OUT8_Mn9@3064_g N_VSS_Mn9@3064_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3065 N_OUT9_Mp9@3065_d N_OUT8_Mp9@3065_g N_VDD_Mp9@3065_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3064 N_OUT9_Mp9@3064_d N_OUT8_Mp9@3064_g N_VDD_Mp9@3064_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3063 N_OUT9_Mn9@3063_d N_OUT8_Mn9@3063_g N_VSS_Mn9@3063_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3062 N_OUT9_Mn9@3062_d N_OUT8_Mn9@3062_g N_VSS_Mn9@3062_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3063 N_OUT9_Mp9@3063_d N_OUT8_Mp9@3063_g N_VDD_Mp9@3063_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3062 N_OUT9_Mp9@3062_d N_OUT8_Mp9@3062_g N_VDD_Mp9@3062_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3061 N_OUT9_Mn9@3061_d N_OUT8_Mn9@3061_g N_VSS_Mn9@3061_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3060 N_OUT9_Mn9@3060_d N_OUT8_Mn9@3060_g N_VSS_Mn9@3060_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3061 N_OUT9_Mp9@3061_d N_OUT8_Mp9@3061_g N_VDD_Mp9@3061_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3060 N_OUT9_Mp9@3060_d N_OUT8_Mp9@3060_g N_VDD_Mp9@3060_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3059 N_OUT9_Mn9@3059_d N_OUT8_Mn9@3059_g N_VSS_Mn9@3059_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3058 N_OUT9_Mn9@3058_d N_OUT8_Mn9@3058_g N_VSS_Mn9@3058_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3059 N_OUT9_Mp9@3059_d N_OUT8_Mp9@3059_g N_VDD_Mp9@3059_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3058 N_OUT9_Mp9@3058_d N_OUT8_Mp9@3058_g N_VDD_Mp9@3058_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3057 N_OUT9_Mn9@3057_d N_OUT8_Mn9@3057_g N_VSS_Mn9@3057_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3056 N_OUT9_Mn9@3056_d N_OUT8_Mn9@3056_g N_VSS_Mn9@3056_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3057 N_OUT9_Mp9@3057_d N_OUT8_Mp9@3057_g N_VDD_Mp9@3057_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3056 N_OUT9_Mp9@3056_d N_OUT8_Mp9@3056_g N_VDD_Mp9@3056_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3055 N_OUT9_Mn9@3055_d N_OUT8_Mn9@3055_g N_VSS_Mn9@3055_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3054 N_OUT9_Mn9@3054_d N_OUT8_Mn9@3054_g N_VSS_Mn9@3054_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3055 N_OUT9_Mp9@3055_d N_OUT8_Mp9@3055_g N_VDD_Mp9@3055_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3054 N_OUT9_Mp9@3054_d N_OUT8_Mp9@3054_g N_VDD_Mp9@3054_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3053 N_OUT9_Mn9@3053_d N_OUT8_Mn9@3053_g N_VSS_Mn9@3053_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3052 N_OUT9_Mn9@3052_d N_OUT8_Mn9@3052_g N_VSS_Mn9@3052_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3053 N_OUT9_Mp9@3053_d N_OUT8_Mp9@3053_g N_VDD_Mp9@3053_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3052 N_OUT9_Mp9@3052_d N_OUT8_Mp9@3052_g N_VDD_Mp9@3052_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3051 N_OUT9_Mn9@3051_d N_OUT8_Mn9@3051_g N_VSS_Mn9@3051_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3050 N_OUT9_Mn9@3050_d N_OUT8_Mn9@3050_g N_VSS_Mn9@3050_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3051 N_OUT9_Mp9@3051_d N_OUT8_Mp9@3051_g N_VDD_Mp9@3051_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3050 N_OUT9_Mp9@3050_d N_OUT8_Mp9@3050_g N_VDD_Mp9@3050_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3049 N_OUT9_Mn9@3049_d N_OUT8_Mn9@3049_g N_VSS_Mn9@3049_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3048 N_OUT9_Mn9@3048_d N_OUT8_Mn9@3048_g N_VSS_Mn9@3048_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3049 N_OUT9_Mp9@3049_d N_OUT8_Mp9@3049_g N_VDD_Mp9@3049_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3048 N_OUT9_Mp9@3048_d N_OUT8_Mp9@3048_g N_VDD_Mp9@3048_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3047 N_OUT9_Mn9@3047_d N_OUT8_Mn9@3047_g N_VSS_Mn9@3047_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3046 N_OUT9_Mn9@3046_d N_OUT8_Mn9@3046_g N_VSS_Mn9@3046_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3047 N_OUT9_Mp9@3047_d N_OUT8_Mp9@3047_g N_VDD_Mp9@3047_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3046 N_OUT9_Mp9@3046_d N_OUT8_Mp9@3046_g N_VDD_Mp9@3046_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3045 N_OUT9_Mn9@3045_d N_OUT8_Mn9@3045_g N_VSS_Mn9@3045_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3044 N_OUT9_Mn9@3044_d N_OUT8_Mn9@3044_g N_VSS_Mn9@3044_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3045 N_OUT9_Mp9@3045_d N_OUT8_Mp9@3045_g N_VDD_Mp9@3045_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3044 N_OUT9_Mp9@3044_d N_OUT8_Mp9@3044_g N_VDD_Mp9@3044_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3043 N_OUT9_Mn9@3043_d N_OUT8_Mn9@3043_g N_VSS_Mn9@3043_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3042 N_OUT9_Mn9@3042_d N_OUT8_Mn9@3042_g N_VSS_Mn9@3042_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3043 N_OUT9_Mp9@3043_d N_OUT8_Mp9@3043_g N_VDD_Mp9@3043_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3042 N_OUT9_Mp9@3042_d N_OUT8_Mp9@3042_g N_VDD_Mp9@3042_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3041 N_OUT9_Mn9@3041_d N_OUT8_Mn9@3041_g N_VSS_Mn9@3041_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3040 N_OUT9_Mn9@3040_d N_OUT8_Mn9@3040_g N_VSS_Mn9@3040_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3041 N_OUT9_Mp9@3041_d N_OUT8_Mp9@3041_g N_VDD_Mp9@3041_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3040 N_OUT9_Mp9@3040_d N_OUT8_Mp9@3040_g N_VDD_Mp9@3040_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3039 N_OUT9_Mn9@3039_d N_OUT8_Mn9@3039_g N_VSS_Mn9@3039_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3038 N_OUT9_Mn9@3038_d N_OUT8_Mn9@3038_g N_VSS_Mn9@3038_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3039 N_OUT9_Mp9@3039_d N_OUT8_Mp9@3039_g N_VDD_Mp9@3039_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3038 N_OUT9_Mp9@3038_d N_OUT8_Mp9@3038_g N_VDD_Mp9@3038_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3037 N_OUT9_Mn9@3037_d N_OUT8_Mn9@3037_g N_VSS_Mn9@3037_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3036 N_OUT9_Mn9@3036_d N_OUT8_Mn9@3036_g N_VSS_Mn9@3036_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3037 N_OUT9_Mp9@3037_d N_OUT8_Mp9@3037_g N_VDD_Mp9@3037_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3036 N_OUT9_Mp9@3036_d N_OUT8_Mp9@3036_g N_VDD_Mp9@3036_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3035 N_OUT9_Mn9@3035_d N_OUT8_Mn9@3035_g N_VSS_Mn9@3035_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3034 N_OUT9_Mn9@3034_d N_OUT8_Mn9@3034_g N_VSS_Mn9@3034_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3035 N_OUT9_Mp9@3035_d N_OUT8_Mp9@3035_g N_VDD_Mp9@3035_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3034 N_OUT9_Mp9@3034_d N_OUT8_Mp9@3034_g N_VDD_Mp9@3034_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3033 N_OUT9_Mn9@3033_d N_OUT8_Mn9@3033_g N_VSS_Mn9@3033_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3032 N_OUT9_Mn9@3032_d N_OUT8_Mn9@3032_g N_VSS_Mn9@3032_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3033 N_OUT9_Mp9@3033_d N_OUT8_Mp9@3033_g N_VDD_Mp9@3033_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3032 N_OUT9_Mp9@3032_d N_OUT8_Mp9@3032_g N_VDD_Mp9@3032_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3031 N_OUT9_Mn9@3031_d N_OUT8_Mn9@3031_g N_VSS_Mn9@3031_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3030 N_OUT9_Mn9@3030_d N_OUT8_Mn9@3030_g N_VSS_Mn9@3030_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3031 N_OUT9_Mp9@3031_d N_OUT8_Mp9@3031_g N_VDD_Mp9@3031_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3030 N_OUT9_Mp9@3030_d N_OUT8_Mp9@3030_g N_VDD_Mp9@3030_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3029 N_OUT9_Mn9@3029_d N_OUT8_Mn9@3029_g N_VSS_Mn9@3029_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3028 N_OUT9_Mn9@3028_d N_OUT8_Mn9@3028_g N_VSS_Mn9@3028_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3029 N_OUT9_Mp9@3029_d N_OUT8_Mp9@3029_g N_VDD_Mp9@3029_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3028 N_OUT9_Mp9@3028_d N_OUT8_Mp9@3028_g N_VDD_Mp9@3028_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3027 N_OUT9_Mn9@3027_d N_OUT8_Mn9@3027_g N_VSS_Mn9@3027_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3026 N_OUT9_Mn9@3026_d N_OUT8_Mn9@3026_g N_VSS_Mn9@3026_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3027 N_OUT9_Mp9@3027_d N_OUT8_Mp9@3027_g N_VDD_Mp9@3027_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3026 N_OUT9_Mp9@3026_d N_OUT8_Mp9@3026_g N_VDD_Mp9@3026_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3025 N_OUT9_Mn9@3025_d N_OUT8_Mn9@3025_g N_VSS_Mn9@3025_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3024 N_OUT9_Mn9@3024_d N_OUT8_Mn9@3024_g N_VSS_Mn9@3024_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3025 N_OUT9_Mp9@3025_d N_OUT8_Mp9@3025_g N_VDD_Mp9@3025_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3024 N_OUT9_Mp9@3024_d N_OUT8_Mp9@3024_g N_VDD_Mp9@3024_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3023 N_OUT9_Mn9@3023_d N_OUT8_Mn9@3023_g N_VSS_Mn9@3023_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3022 N_OUT9_Mn9@3022_d N_OUT8_Mn9@3022_g N_VSS_Mn9@3022_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3023 N_OUT9_Mp9@3023_d N_OUT8_Mp9@3023_g N_VDD_Mp9@3023_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3022 N_OUT9_Mp9@3022_d N_OUT8_Mp9@3022_g N_VDD_Mp9@3022_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3021 N_OUT9_Mn9@3021_d N_OUT8_Mn9@3021_g N_VSS_Mn9@3021_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3020 N_OUT9_Mn9@3020_d N_OUT8_Mn9@3020_g N_VSS_Mn9@3020_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3021 N_OUT9_Mp9@3021_d N_OUT8_Mp9@3021_g N_VDD_Mp9@3021_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3020 N_OUT9_Mp9@3020_d N_OUT8_Mp9@3020_g N_VDD_Mp9@3020_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3019 N_OUT9_Mn9@3019_d N_OUT8_Mn9@3019_g N_VSS_Mn9@3019_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3018 N_OUT9_Mn9@3018_d N_OUT8_Mn9@3018_g N_VSS_Mn9@3018_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3019 N_OUT9_Mp9@3019_d N_OUT8_Mp9@3019_g N_VDD_Mp9@3019_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3018 N_OUT9_Mp9@3018_d N_OUT8_Mp9@3018_g N_VDD_Mp9@3018_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3017 N_OUT9_Mn9@3017_d N_OUT8_Mn9@3017_g N_VSS_Mn9@3017_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3016 N_OUT9_Mn9@3016_d N_OUT8_Mn9@3016_g N_VSS_Mn9@3016_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3017 N_OUT9_Mp9@3017_d N_OUT8_Mp9@3017_g N_VDD_Mp9@3017_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3016 N_OUT9_Mp9@3016_d N_OUT8_Mp9@3016_g N_VDD_Mp9@3016_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3015 N_OUT9_Mn9@3015_d N_OUT8_Mn9@3015_g N_VSS_Mn9@3015_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3014 N_OUT9_Mn9@3014_d N_OUT8_Mn9@3014_g N_VSS_Mn9@3014_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3015 N_OUT9_Mp9@3015_d N_OUT8_Mp9@3015_g N_VDD_Mp9@3015_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3014 N_OUT9_Mp9@3014_d N_OUT8_Mp9@3014_g N_VDD_Mp9@3014_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3013 N_OUT9_Mn9@3013_d N_OUT8_Mn9@3013_g N_VSS_Mn9@3013_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3012 N_OUT9_Mn9@3012_d N_OUT8_Mn9@3012_g N_VSS_Mn9@3012_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3013 N_OUT9_Mp9@3013_d N_OUT8_Mp9@3013_g N_VDD_Mp9@3013_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3012 N_OUT9_Mp9@3012_d N_OUT8_Mp9@3012_g N_VDD_Mp9@3012_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3011 N_OUT9_Mn9@3011_d N_OUT8_Mn9@3011_g N_VSS_Mn9@3011_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3010 N_OUT9_Mn9@3010_d N_OUT8_Mn9@3010_g N_VSS_Mn9@3010_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3011 N_OUT9_Mp9@3011_d N_OUT8_Mp9@3011_g N_VDD_Mp9@3011_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3010 N_OUT9_Mp9@3010_d N_OUT8_Mp9@3010_g N_VDD_Mp9@3010_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3009 N_OUT9_Mn9@3009_d N_OUT8_Mn9@3009_g N_VSS_Mn9@3009_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3008 N_OUT9_Mn9@3008_d N_OUT8_Mn9@3008_g N_VSS_Mn9@3008_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3009 N_OUT9_Mp9@3009_d N_OUT8_Mp9@3009_g N_VDD_Mp9@3009_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3008 N_OUT9_Mp9@3008_d N_OUT8_Mp9@3008_g N_VDD_Mp9@3008_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3007 N_OUT9_Mn9@3007_d N_OUT8_Mn9@3007_g N_VSS_Mn9@3007_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3006 N_OUT9_Mn9@3006_d N_OUT8_Mn9@3006_g N_VSS_Mn9@3006_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3007 N_OUT9_Mp9@3007_d N_OUT8_Mp9@3007_g N_VDD_Mp9@3007_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3006 N_OUT9_Mp9@3006_d N_OUT8_Mp9@3006_g N_VDD_Mp9@3006_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3005 N_OUT9_Mn9@3005_d N_OUT8_Mn9@3005_g N_VSS_Mn9@3005_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3004 N_OUT9_Mn9@3004_d N_OUT8_Mn9@3004_g N_VSS_Mn9@3004_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3005 N_OUT9_Mp9@3005_d N_OUT8_Mp9@3005_g N_VDD_Mp9@3005_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3004 N_OUT9_Mp9@3004_d N_OUT8_Mp9@3004_g N_VDD_Mp9@3004_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3003 N_OUT9_Mn9@3003_d N_OUT8_Mn9@3003_g N_VSS_Mn9@3003_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3002 N_OUT9_Mn9@3002_d N_OUT8_Mn9@3002_g N_VSS_Mn9@3002_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3003 N_OUT9_Mp9@3003_d N_OUT8_Mp9@3003_g N_VDD_Mp9@3003_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3002 N_OUT9_Mp9@3002_d N_OUT8_Mp9@3002_g N_VDD_Mp9@3002_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3001 N_OUT9_Mn9@3001_d N_OUT8_Mn9@3001_g N_VSS_Mn9@3001_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@3000 N_OUT9_Mn9@3000_d N_OUT8_Mn9@3000_g N_VSS_Mn9@3000_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3001 N_OUT9_Mp9@3001_d N_OUT8_Mp9@3001_g N_VDD_Mp9@3001_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@3000 N_OUT9_Mp9@3000_d N_OUT8_Mp9@3000_g N_VDD_Mp9@3000_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2999 N_OUT9_Mn9@2999_d N_OUT8_Mn9@2999_g N_VSS_Mn9@2999_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2998 N_OUT9_Mn9@2998_d N_OUT8_Mn9@2998_g N_VSS_Mn9@2998_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2999 N_OUT9_Mp9@2999_d N_OUT8_Mp9@2999_g N_VDD_Mp9@2999_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2998 N_OUT9_Mp9@2998_d N_OUT8_Mp9@2998_g N_VDD_Mp9@2998_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2997 N_OUT9_Mn9@2997_d N_OUT8_Mn9@2997_g N_VSS_Mn9@2997_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2996 N_OUT9_Mn9@2996_d N_OUT8_Mn9@2996_g N_VSS_Mn9@2996_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2997 N_OUT9_Mp9@2997_d N_OUT8_Mp9@2997_g N_VDD_Mp9@2997_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2996 N_OUT9_Mp9@2996_d N_OUT8_Mp9@2996_g N_VDD_Mp9@2996_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2995 N_OUT9_Mn9@2995_d N_OUT8_Mn9@2995_g N_VSS_Mn9@2995_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2994 N_OUT9_Mn9@2994_d N_OUT8_Mn9@2994_g N_VSS_Mn9@2994_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2995 N_OUT9_Mp9@2995_d N_OUT8_Mp9@2995_g N_VDD_Mp9@2995_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2994 N_OUT9_Mp9@2994_d N_OUT8_Mp9@2994_g N_VDD_Mp9@2994_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2993 N_OUT9_Mn9@2993_d N_OUT8_Mn9@2993_g N_VSS_Mn9@2993_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2992 N_OUT9_Mn9@2992_d N_OUT8_Mn9@2992_g N_VSS_Mn9@2992_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2993 N_OUT9_Mp9@2993_d N_OUT8_Mp9@2993_g N_VDD_Mp9@2993_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2992 N_OUT9_Mp9@2992_d N_OUT8_Mp9@2992_g N_VDD_Mp9@2992_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2991 N_OUT9_Mn9@2991_d N_OUT8_Mn9@2991_g N_VSS_Mn9@2991_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2990 N_OUT9_Mn9@2990_d N_OUT8_Mn9@2990_g N_VSS_Mn9@2990_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2991 N_OUT9_Mp9@2991_d N_OUT8_Mp9@2991_g N_VDD_Mp9@2991_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2990 N_OUT9_Mp9@2990_d N_OUT8_Mp9@2990_g N_VDD_Mp9@2990_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2989 N_OUT9_Mn9@2989_d N_OUT8_Mn9@2989_g N_VSS_Mn9@2989_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2988 N_OUT9_Mn9@2988_d N_OUT8_Mn9@2988_g N_VSS_Mn9@2988_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2989 N_OUT9_Mp9@2989_d N_OUT8_Mp9@2989_g N_VDD_Mp9@2989_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2988 N_OUT9_Mp9@2988_d N_OUT8_Mp9@2988_g N_VDD_Mp9@2988_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2987 N_OUT9_Mn9@2987_d N_OUT8_Mn9@2987_g N_VSS_Mn9@2987_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2986 N_OUT9_Mn9@2986_d N_OUT8_Mn9@2986_g N_VSS_Mn9@2986_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2987 N_OUT9_Mp9@2987_d N_OUT8_Mp9@2987_g N_VDD_Mp9@2987_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2986 N_OUT9_Mp9@2986_d N_OUT8_Mp9@2986_g N_VDD_Mp9@2986_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2985 N_OUT9_Mn9@2985_d N_OUT8_Mn9@2985_g N_VSS_Mn9@2985_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2984 N_OUT9_Mn9@2984_d N_OUT8_Mn9@2984_g N_VSS_Mn9@2984_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2985 N_OUT9_Mp9@2985_d N_OUT8_Mp9@2985_g N_VDD_Mp9@2985_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2984 N_OUT9_Mp9@2984_d N_OUT8_Mp9@2984_g N_VDD_Mp9@2984_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2983 N_OUT9_Mn9@2983_d N_OUT8_Mn9@2983_g N_VSS_Mn9@2983_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2982 N_OUT9_Mn9@2982_d N_OUT8_Mn9@2982_g N_VSS_Mn9@2982_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2983 N_OUT9_Mp9@2983_d N_OUT8_Mp9@2983_g N_VDD_Mp9@2983_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2982 N_OUT9_Mp9@2982_d N_OUT8_Mp9@2982_g N_VDD_Mp9@2982_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2981 N_OUT9_Mn9@2981_d N_OUT8_Mn9@2981_g N_VSS_Mn9@2981_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2980 N_OUT9_Mn9@2980_d N_OUT8_Mn9@2980_g N_VSS_Mn9@2980_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2981 N_OUT9_Mp9@2981_d N_OUT8_Mp9@2981_g N_VDD_Mp9@2981_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2980 N_OUT9_Mp9@2980_d N_OUT8_Mp9@2980_g N_VDD_Mp9@2980_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2979 N_OUT9_Mn9@2979_d N_OUT8_Mn9@2979_g N_VSS_Mn9@2979_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2978 N_OUT9_Mn9@2978_d N_OUT8_Mn9@2978_g N_VSS_Mn9@2978_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2979 N_OUT9_Mp9@2979_d N_OUT8_Mp9@2979_g N_VDD_Mp9@2979_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2978 N_OUT9_Mp9@2978_d N_OUT8_Mp9@2978_g N_VDD_Mp9@2978_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2977 N_OUT9_Mn9@2977_d N_OUT8_Mn9@2977_g N_VSS_Mn9@2977_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2976 N_OUT9_Mn9@2976_d N_OUT8_Mn9@2976_g N_VSS_Mn9@2976_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2977 N_OUT9_Mp9@2977_d N_OUT8_Mp9@2977_g N_VDD_Mp9@2977_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2976 N_OUT9_Mp9@2976_d N_OUT8_Mp9@2976_g N_VDD_Mp9@2976_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2975 N_OUT9_Mn9@2975_d N_OUT8_Mn9@2975_g N_VSS_Mn9@2975_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2974 N_OUT9_Mn9@2974_d N_OUT8_Mn9@2974_g N_VSS_Mn9@2974_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2975 N_OUT9_Mp9@2975_d N_OUT8_Mp9@2975_g N_VDD_Mp9@2975_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2974 N_OUT9_Mp9@2974_d N_OUT8_Mp9@2974_g N_VDD_Mp9@2974_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2973 N_OUT9_Mn9@2973_d N_OUT8_Mn9@2973_g N_VSS_Mn9@2973_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2972 N_OUT9_Mn9@2972_d N_OUT8_Mn9@2972_g N_VSS_Mn9@2972_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2973 N_OUT9_Mp9@2973_d N_OUT8_Mp9@2973_g N_VDD_Mp9@2973_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2972 N_OUT9_Mp9@2972_d N_OUT8_Mp9@2972_g N_VDD_Mp9@2972_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2971 N_OUT9_Mn9@2971_d N_OUT8_Mn9@2971_g N_VSS_Mn9@2971_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2970 N_OUT9_Mn9@2970_d N_OUT8_Mn9@2970_g N_VSS_Mn9@2970_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2971 N_OUT9_Mp9@2971_d N_OUT8_Mp9@2971_g N_VDD_Mp9@2971_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2970 N_OUT9_Mp9@2970_d N_OUT8_Mp9@2970_g N_VDD_Mp9@2970_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2969 N_OUT9_Mn9@2969_d N_OUT8_Mn9@2969_g N_VSS_Mn9@2969_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2968 N_OUT9_Mn9@2968_d N_OUT8_Mn9@2968_g N_VSS_Mn9@2968_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2969 N_OUT9_Mp9@2969_d N_OUT8_Mp9@2969_g N_VDD_Mp9@2969_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2968 N_OUT9_Mp9@2968_d N_OUT8_Mp9@2968_g N_VDD_Mp9@2968_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2967 N_OUT9_Mn9@2967_d N_OUT8_Mn9@2967_g N_VSS_Mn9@2967_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2966 N_OUT9_Mn9@2966_d N_OUT8_Mn9@2966_g N_VSS_Mn9@2966_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2967 N_OUT9_Mp9@2967_d N_OUT8_Mp9@2967_g N_VDD_Mp9@2967_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2966 N_OUT9_Mp9@2966_d N_OUT8_Mp9@2966_g N_VDD_Mp9@2966_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2965 N_OUT9_Mn9@2965_d N_OUT8_Mn9@2965_g N_VSS_Mn9@2965_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2964 N_OUT9_Mn9@2964_d N_OUT8_Mn9@2964_g N_VSS_Mn9@2964_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2965 N_OUT9_Mp9@2965_d N_OUT8_Mp9@2965_g N_VDD_Mp9@2965_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2964 N_OUT9_Mp9@2964_d N_OUT8_Mp9@2964_g N_VDD_Mp9@2964_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2963 N_OUT9_Mn9@2963_d N_OUT8_Mn9@2963_g N_VSS_Mn9@2963_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2962 N_OUT9_Mn9@2962_d N_OUT8_Mn9@2962_g N_VSS_Mn9@2962_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2963 N_OUT9_Mp9@2963_d N_OUT8_Mp9@2963_g N_VDD_Mp9@2963_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2962 N_OUT9_Mp9@2962_d N_OUT8_Mp9@2962_g N_VDD_Mp9@2962_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2961 N_OUT9_Mn9@2961_d N_OUT8_Mn9@2961_g N_VSS_Mn9@2961_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2960 N_OUT9_Mn9@2960_d N_OUT8_Mn9@2960_g N_VSS_Mn9@2960_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2961 N_OUT9_Mp9@2961_d N_OUT8_Mp9@2961_g N_VDD_Mp9@2961_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2960 N_OUT9_Mp9@2960_d N_OUT8_Mp9@2960_g N_VDD_Mp9@2960_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2959 N_OUT9_Mn9@2959_d N_OUT8_Mn9@2959_g N_VSS_Mn9@2959_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2958 N_OUT9_Mn9@2958_d N_OUT8_Mn9@2958_g N_VSS_Mn9@2958_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2959 N_OUT9_Mp9@2959_d N_OUT8_Mp9@2959_g N_VDD_Mp9@2959_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2958 N_OUT9_Mp9@2958_d N_OUT8_Mp9@2958_g N_VDD_Mp9@2958_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2957 N_OUT9_Mn9@2957_d N_OUT8_Mn9@2957_g N_VSS_Mn9@2957_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2956 N_OUT9_Mn9@2956_d N_OUT8_Mn9@2956_g N_VSS_Mn9@2956_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2957 N_OUT9_Mp9@2957_d N_OUT8_Mp9@2957_g N_VDD_Mp9@2957_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2956 N_OUT9_Mp9@2956_d N_OUT8_Mp9@2956_g N_VDD_Mp9@2956_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2955 N_OUT9_Mn9@2955_d N_OUT8_Mn9@2955_g N_VSS_Mn9@2955_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2954 N_OUT9_Mn9@2954_d N_OUT8_Mn9@2954_g N_VSS_Mn9@2954_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2955 N_OUT9_Mp9@2955_d N_OUT8_Mp9@2955_g N_VDD_Mp9@2955_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2954 N_OUT9_Mp9@2954_d N_OUT8_Mp9@2954_g N_VDD_Mp9@2954_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2953 N_OUT9_Mn9@2953_d N_OUT8_Mn9@2953_g N_VSS_Mn9@2953_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2952 N_OUT9_Mn9@2952_d N_OUT8_Mn9@2952_g N_VSS_Mn9@2952_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2953 N_OUT9_Mp9@2953_d N_OUT8_Mp9@2953_g N_VDD_Mp9@2953_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2952 N_OUT9_Mp9@2952_d N_OUT8_Mp9@2952_g N_VDD_Mp9@2952_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2951 N_OUT9_Mn9@2951_d N_OUT8_Mn9@2951_g N_VSS_Mn9@2951_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2950 N_OUT9_Mn9@2950_d N_OUT8_Mn9@2950_g N_VSS_Mn9@2950_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2951 N_OUT9_Mp9@2951_d N_OUT8_Mp9@2951_g N_VDD_Mp9@2951_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2950 N_OUT9_Mp9@2950_d N_OUT8_Mp9@2950_g N_VDD_Mp9@2950_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2949 N_OUT9_Mn9@2949_d N_OUT8_Mn9@2949_g N_VSS_Mn9@2949_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2948 N_OUT9_Mn9@2948_d N_OUT8_Mn9@2948_g N_VSS_Mn9@2948_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2949 N_OUT9_Mp9@2949_d N_OUT8_Mp9@2949_g N_VDD_Mp9@2949_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2948 N_OUT9_Mp9@2948_d N_OUT8_Mp9@2948_g N_VDD_Mp9@2948_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2947 N_OUT9_Mn9@2947_d N_OUT8_Mn9@2947_g N_VSS_Mn9@2947_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2946 N_OUT9_Mn9@2946_d N_OUT8_Mn9@2946_g N_VSS_Mn9@2946_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2947 N_OUT9_Mp9@2947_d N_OUT8_Mp9@2947_g N_VDD_Mp9@2947_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2946 N_OUT9_Mp9@2946_d N_OUT8_Mp9@2946_g N_VDD_Mp9@2946_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2945 N_OUT9_Mn9@2945_d N_OUT8_Mn9@2945_g N_VSS_Mn9@2945_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2944 N_OUT9_Mn9@2944_d N_OUT8_Mn9@2944_g N_VSS_Mn9@2944_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2945 N_OUT9_Mp9@2945_d N_OUT8_Mp9@2945_g N_VDD_Mp9@2945_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2944 N_OUT9_Mp9@2944_d N_OUT8_Mp9@2944_g N_VDD_Mp9@2944_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2943 N_OUT9_Mn9@2943_d N_OUT8_Mn9@2943_g N_VSS_Mn9@2943_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2942 N_OUT9_Mn9@2942_d N_OUT8_Mn9@2942_g N_VSS_Mn9@2942_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2943 N_OUT9_Mp9@2943_d N_OUT8_Mp9@2943_g N_VDD_Mp9@2943_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2942 N_OUT9_Mp9@2942_d N_OUT8_Mp9@2942_g N_VDD_Mp9@2942_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2941 N_OUT9_Mn9@2941_d N_OUT8_Mn9@2941_g N_VSS_Mn9@2941_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2940 N_OUT9_Mn9@2940_d N_OUT8_Mn9@2940_g N_VSS_Mn9@2940_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2941 N_OUT9_Mp9@2941_d N_OUT8_Mp9@2941_g N_VDD_Mp9@2941_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2940 N_OUT9_Mp9@2940_d N_OUT8_Mp9@2940_g N_VDD_Mp9@2940_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2939 N_OUT9_Mn9@2939_d N_OUT8_Mn9@2939_g N_VSS_Mn9@2939_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2938 N_OUT9_Mn9@2938_d N_OUT8_Mn9@2938_g N_VSS_Mn9@2938_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2939 N_OUT9_Mp9@2939_d N_OUT8_Mp9@2939_g N_VDD_Mp9@2939_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2938 N_OUT9_Mp9@2938_d N_OUT8_Mp9@2938_g N_VDD_Mp9@2938_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2937 N_OUT9_Mn9@2937_d N_OUT8_Mn9@2937_g N_VSS_Mn9@2937_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2936 N_OUT9_Mn9@2936_d N_OUT8_Mn9@2936_g N_VSS_Mn9@2936_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2937 N_OUT9_Mp9@2937_d N_OUT8_Mp9@2937_g N_VDD_Mp9@2937_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2936 N_OUT9_Mp9@2936_d N_OUT8_Mp9@2936_g N_VDD_Mp9@2936_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2935 N_OUT9_Mn9@2935_d N_OUT8_Mn9@2935_g N_VSS_Mn9@2935_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2934 N_OUT9_Mn9@2934_d N_OUT8_Mn9@2934_g N_VSS_Mn9@2934_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2935 N_OUT9_Mp9@2935_d N_OUT8_Mp9@2935_g N_VDD_Mp9@2935_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2934 N_OUT9_Mp9@2934_d N_OUT8_Mp9@2934_g N_VDD_Mp9@2934_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2933 N_OUT9_Mn9@2933_d N_OUT8_Mn9@2933_g N_VSS_Mn9@2933_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2932 N_OUT9_Mn9@2932_d N_OUT8_Mn9@2932_g N_VSS_Mn9@2932_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2933 N_OUT9_Mp9@2933_d N_OUT8_Mp9@2933_g N_VDD_Mp9@2933_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2932 N_OUT9_Mp9@2932_d N_OUT8_Mp9@2932_g N_VDD_Mp9@2932_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2931 N_OUT9_Mn9@2931_d N_OUT8_Mn9@2931_g N_VSS_Mn9@2931_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2930 N_OUT9_Mn9@2930_d N_OUT8_Mn9@2930_g N_VSS_Mn9@2930_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2931 N_OUT9_Mp9@2931_d N_OUT8_Mp9@2931_g N_VDD_Mp9@2931_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2930 N_OUT9_Mp9@2930_d N_OUT8_Mp9@2930_g N_VDD_Mp9@2930_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2929 N_OUT9_Mn9@2929_d N_OUT8_Mn9@2929_g N_VSS_Mn9@2929_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2928 N_OUT9_Mn9@2928_d N_OUT8_Mn9@2928_g N_VSS_Mn9@2928_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2929 N_OUT9_Mp9@2929_d N_OUT8_Mp9@2929_g N_VDD_Mp9@2929_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2928 N_OUT9_Mp9@2928_d N_OUT8_Mp9@2928_g N_VDD_Mp9@2928_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2927 N_OUT9_Mn9@2927_d N_OUT8_Mn9@2927_g N_VSS_Mn9@2927_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2926 N_OUT9_Mn9@2926_d N_OUT8_Mn9@2926_g N_VSS_Mn9@2926_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2927 N_OUT9_Mp9@2927_d N_OUT8_Mp9@2927_g N_VDD_Mp9@2927_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2926 N_OUT9_Mp9@2926_d N_OUT8_Mp9@2926_g N_VDD_Mp9@2926_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2925 N_OUT9_Mn9@2925_d N_OUT8_Mn9@2925_g N_VSS_Mn9@2925_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2924 N_OUT9_Mn9@2924_d N_OUT8_Mn9@2924_g N_VSS_Mn9@2924_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2925 N_OUT9_Mp9@2925_d N_OUT8_Mp9@2925_g N_VDD_Mp9@2925_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2924 N_OUT9_Mp9@2924_d N_OUT8_Mp9@2924_g N_VDD_Mp9@2924_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2923 N_OUT9_Mn9@2923_d N_OUT8_Mn9@2923_g N_VSS_Mn9@2923_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2922 N_OUT9_Mn9@2922_d N_OUT8_Mn9@2922_g N_VSS_Mn9@2922_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2923 N_OUT9_Mp9@2923_d N_OUT8_Mp9@2923_g N_VDD_Mp9@2923_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2922 N_OUT9_Mp9@2922_d N_OUT8_Mp9@2922_g N_VDD_Mp9@2922_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2921 N_OUT9_Mn9@2921_d N_OUT8_Mn9@2921_g N_VSS_Mn9@2921_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2920 N_OUT9_Mn9@2920_d N_OUT8_Mn9@2920_g N_VSS_Mn9@2920_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2921 N_OUT9_Mp9@2921_d N_OUT8_Mp9@2921_g N_VDD_Mp9@2921_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2920 N_OUT9_Mp9@2920_d N_OUT8_Mp9@2920_g N_VDD_Mp9@2920_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2919 N_OUT9_Mn9@2919_d N_OUT8_Mn9@2919_g N_VSS_Mn9@2919_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2918 N_OUT9_Mn9@2918_d N_OUT8_Mn9@2918_g N_VSS_Mn9@2918_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2919 N_OUT9_Mp9@2919_d N_OUT8_Mp9@2919_g N_VDD_Mp9@2919_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2918 N_OUT9_Mp9@2918_d N_OUT8_Mp9@2918_g N_VDD_Mp9@2918_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2917 N_OUT9_Mn9@2917_d N_OUT8_Mn9@2917_g N_VSS_Mn9@2917_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2916 N_OUT9_Mn9@2916_d N_OUT8_Mn9@2916_g N_VSS_Mn9@2916_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2917 N_OUT9_Mp9@2917_d N_OUT8_Mp9@2917_g N_VDD_Mp9@2917_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2916 N_OUT9_Mp9@2916_d N_OUT8_Mp9@2916_g N_VDD_Mp9@2916_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2915 N_OUT9_Mn9@2915_d N_OUT8_Mn9@2915_g N_VSS_Mn9@2915_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2914 N_OUT9_Mn9@2914_d N_OUT8_Mn9@2914_g N_VSS_Mn9@2914_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2915 N_OUT9_Mp9@2915_d N_OUT8_Mp9@2915_g N_VDD_Mp9@2915_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2914 N_OUT9_Mp9@2914_d N_OUT8_Mp9@2914_g N_VDD_Mp9@2914_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2913 N_OUT9_Mn9@2913_d N_OUT8_Mn9@2913_g N_VSS_Mn9@2913_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2912 N_OUT9_Mn9@2912_d N_OUT8_Mn9@2912_g N_VSS_Mn9@2912_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2913 N_OUT9_Mp9@2913_d N_OUT8_Mp9@2913_g N_VDD_Mp9@2913_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2912 N_OUT9_Mp9@2912_d N_OUT8_Mp9@2912_g N_VDD_Mp9@2912_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2911 N_OUT9_Mn9@2911_d N_OUT8_Mn9@2911_g N_VSS_Mn9@2911_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2910 N_OUT9_Mn9@2910_d N_OUT8_Mn9@2910_g N_VSS_Mn9@2910_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2911 N_OUT9_Mp9@2911_d N_OUT8_Mp9@2911_g N_VDD_Mp9@2911_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2910 N_OUT9_Mp9@2910_d N_OUT8_Mp9@2910_g N_VDD_Mp9@2910_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2909 N_OUT9_Mn9@2909_d N_OUT8_Mn9@2909_g N_VSS_Mn9@2909_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2908 N_OUT9_Mn9@2908_d N_OUT8_Mn9@2908_g N_VSS_Mn9@2908_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2909 N_OUT9_Mp9@2909_d N_OUT8_Mp9@2909_g N_VDD_Mp9@2909_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2908 N_OUT9_Mp9@2908_d N_OUT8_Mp9@2908_g N_VDD_Mp9@2908_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2907 N_OUT9_Mn9@2907_d N_OUT8_Mn9@2907_g N_VSS_Mn9@2907_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2906 N_OUT9_Mn9@2906_d N_OUT8_Mn9@2906_g N_VSS_Mn9@2906_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2907 N_OUT9_Mp9@2907_d N_OUT8_Mp9@2907_g N_VDD_Mp9@2907_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2906 N_OUT9_Mp9@2906_d N_OUT8_Mp9@2906_g N_VDD_Mp9@2906_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2905 N_OUT9_Mn9@2905_d N_OUT8_Mn9@2905_g N_VSS_Mn9@2905_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2904 N_OUT9_Mn9@2904_d N_OUT8_Mn9@2904_g N_VSS_Mn9@2904_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2905 N_OUT9_Mp9@2905_d N_OUT8_Mp9@2905_g N_VDD_Mp9@2905_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2904 N_OUT9_Mp9@2904_d N_OUT8_Mp9@2904_g N_VDD_Mp9@2904_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2903 N_OUT9_Mn9@2903_d N_OUT8_Mn9@2903_g N_VSS_Mn9@2903_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2902 N_OUT9_Mn9@2902_d N_OUT8_Mn9@2902_g N_VSS_Mn9@2902_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2903 N_OUT9_Mp9@2903_d N_OUT8_Mp9@2903_g N_VDD_Mp9@2903_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2902 N_OUT9_Mp9@2902_d N_OUT8_Mp9@2902_g N_VDD_Mp9@2902_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2901 N_OUT9_Mn9@2901_d N_OUT8_Mn9@2901_g N_VSS_Mn9@2901_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2900 N_OUT9_Mn9@2900_d N_OUT8_Mn9@2900_g N_VSS_Mn9@2900_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2901 N_OUT9_Mp9@2901_d N_OUT8_Mp9@2901_g N_VDD_Mp9@2901_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2900 N_OUT9_Mp9@2900_d N_OUT8_Mp9@2900_g N_VDD_Mp9@2900_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2899 N_OUT9_Mn9@2899_d N_OUT8_Mn9@2899_g N_VSS_Mn9@2899_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2898 N_OUT9_Mn9@2898_d N_OUT8_Mn9@2898_g N_VSS_Mn9@2898_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2899 N_OUT9_Mp9@2899_d N_OUT8_Mp9@2899_g N_VDD_Mp9@2899_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2898 N_OUT9_Mp9@2898_d N_OUT8_Mp9@2898_g N_VDD_Mp9@2898_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2897 N_OUT9_Mn9@2897_d N_OUT8_Mn9@2897_g N_VSS_Mn9@2897_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2896 N_OUT9_Mn9@2896_d N_OUT8_Mn9@2896_g N_VSS_Mn9@2896_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2897 N_OUT9_Mp9@2897_d N_OUT8_Mp9@2897_g N_VDD_Mp9@2897_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2896 N_OUT9_Mp9@2896_d N_OUT8_Mp9@2896_g N_VDD_Mp9@2896_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2895 N_OUT9_Mn9@2895_d N_OUT8_Mn9@2895_g N_VSS_Mn9@2895_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2894 N_OUT9_Mn9@2894_d N_OUT8_Mn9@2894_g N_VSS_Mn9@2894_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2895 N_OUT9_Mp9@2895_d N_OUT8_Mp9@2895_g N_VDD_Mp9@2895_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2894 N_OUT9_Mp9@2894_d N_OUT8_Mp9@2894_g N_VDD_Mp9@2894_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2893 N_OUT9_Mn9@2893_d N_OUT8_Mn9@2893_g N_VSS_Mn9@2893_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2892 N_OUT9_Mn9@2892_d N_OUT8_Mn9@2892_g N_VSS_Mn9@2892_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2893 N_OUT9_Mp9@2893_d N_OUT8_Mp9@2893_g N_VDD_Mp9@2893_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2892 N_OUT9_Mp9@2892_d N_OUT8_Mp9@2892_g N_VDD_Mp9@2892_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2891 N_OUT9_Mn9@2891_d N_OUT8_Mn9@2891_g N_VSS_Mn9@2891_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2890 N_OUT9_Mn9@2890_d N_OUT8_Mn9@2890_g N_VSS_Mn9@2890_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2891 N_OUT9_Mp9@2891_d N_OUT8_Mp9@2891_g N_VDD_Mp9@2891_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2890 N_OUT9_Mp9@2890_d N_OUT8_Mp9@2890_g N_VDD_Mp9@2890_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2889 N_OUT9_Mn9@2889_d N_OUT8_Mn9@2889_g N_VSS_Mn9@2889_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2888 N_OUT9_Mn9@2888_d N_OUT8_Mn9@2888_g N_VSS_Mn9@2888_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2889 N_OUT9_Mp9@2889_d N_OUT8_Mp9@2889_g N_VDD_Mp9@2889_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2888 N_OUT9_Mp9@2888_d N_OUT8_Mp9@2888_g N_VDD_Mp9@2888_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2887 N_OUT9_Mn9@2887_d N_OUT8_Mn9@2887_g N_VSS_Mn9@2887_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2886 N_OUT9_Mn9@2886_d N_OUT8_Mn9@2886_g N_VSS_Mn9@2886_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2887 N_OUT9_Mp9@2887_d N_OUT8_Mp9@2887_g N_VDD_Mp9@2887_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2886 N_OUT9_Mp9@2886_d N_OUT8_Mp9@2886_g N_VDD_Mp9@2886_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2885 N_OUT9_Mn9@2885_d N_OUT8_Mn9@2885_g N_VSS_Mn9@2885_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2884 N_OUT9_Mn9@2884_d N_OUT8_Mn9@2884_g N_VSS_Mn9@2884_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2885 N_OUT9_Mp9@2885_d N_OUT8_Mp9@2885_g N_VDD_Mp9@2885_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2884 N_OUT9_Mp9@2884_d N_OUT8_Mp9@2884_g N_VDD_Mp9@2884_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2883 N_OUT9_Mn9@2883_d N_OUT8_Mn9@2883_g N_VSS_Mn9@2883_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2882 N_OUT9_Mn9@2882_d N_OUT8_Mn9@2882_g N_VSS_Mn9@2882_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2883 N_OUT9_Mp9@2883_d N_OUT8_Mp9@2883_g N_VDD_Mp9@2883_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2882 N_OUT9_Mp9@2882_d N_OUT8_Mp9@2882_g N_VDD_Mp9@2882_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2881 N_OUT9_Mn9@2881_d N_OUT8_Mn9@2881_g N_VSS_Mn9@2881_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2880 N_OUT9_Mn9@2880_d N_OUT8_Mn9@2880_g N_VSS_Mn9@2880_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2881 N_OUT9_Mp9@2881_d N_OUT8_Mp9@2881_g N_VDD_Mp9@2881_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2880 N_OUT9_Mp9@2880_d N_OUT8_Mp9@2880_g N_VDD_Mp9@2880_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2879 N_OUT9_Mn9@2879_d N_OUT8_Mn9@2879_g N_VSS_Mn9@2879_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2878 N_OUT9_Mn9@2878_d N_OUT8_Mn9@2878_g N_VSS_Mn9@2878_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2879 N_OUT9_Mp9@2879_d N_OUT8_Mp9@2879_g N_VDD_Mp9@2879_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2878 N_OUT9_Mp9@2878_d N_OUT8_Mp9@2878_g N_VDD_Mp9@2878_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2877 N_OUT9_Mn9@2877_d N_OUT8_Mn9@2877_g N_VSS_Mn9@2877_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2876 N_OUT9_Mn9@2876_d N_OUT8_Mn9@2876_g N_VSS_Mn9@2876_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2877 N_OUT9_Mp9@2877_d N_OUT8_Mp9@2877_g N_VDD_Mp9@2877_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2876 N_OUT9_Mp9@2876_d N_OUT8_Mp9@2876_g N_VDD_Mp9@2876_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2875 N_OUT9_Mn9@2875_d N_OUT8_Mn9@2875_g N_VSS_Mn9@2875_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2874 N_OUT9_Mn9@2874_d N_OUT8_Mn9@2874_g N_VSS_Mn9@2874_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2875 N_OUT9_Mp9@2875_d N_OUT8_Mp9@2875_g N_VDD_Mp9@2875_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2874 N_OUT9_Mp9@2874_d N_OUT8_Mp9@2874_g N_VDD_Mp9@2874_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2873 N_OUT9_Mn9@2873_d N_OUT8_Mn9@2873_g N_VSS_Mn9@2873_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2872 N_OUT9_Mn9@2872_d N_OUT8_Mn9@2872_g N_VSS_Mn9@2872_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2873 N_OUT9_Mp9@2873_d N_OUT8_Mp9@2873_g N_VDD_Mp9@2873_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2872 N_OUT9_Mp9@2872_d N_OUT8_Mp9@2872_g N_VDD_Mp9@2872_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2871 N_OUT9_Mn9@2871_d N_OUT8_Mn9@2871_g N_VSS_Mn9@2871_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2870 N_OUT9_Mn9@2870_d N_OUT8_Mn9@2870_g N_VSS_Mn9@2870_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2871 N_OUT9_Mp9@2871_d N_OUT8_Mp9@2871_g N_VDD_Mp9@2871_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2870 N_OUT9_Mp9@2870_d N_OUT8_Mp9@2870_g N_VDD_Mp9@2870_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2869 N_OUT9_Mn9@2869_d N_OUT8_Mn9@2869_g N_VSS_Mn9@2869_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2868 N_OUT9_Mn9@2868_d N_OUT8_Mn9@2868_g N_VSS_Mn9@2868_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2869 N_OUT9_Mp9@2869_d N_OUT8_Mp9@2869_g N_VDD_Mp9@2869_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2868 N_OUT9_Mp9@2868_d N_OUT8_Mp9@2868_g N_VDD_Mp9@2868_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2867 N_OUT9_Mn9@2867_d N_OUT8_Mn9@2867_g N_VSS_Mn9@2867_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2866 N_OUT9_Mn9@2866_d N_OUT8_Mn9@2866_g N_VSS_Mn9@2866_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2867 N_OUT9_Mp9@2867_d N_OUT8_Mp9@2867_g N_VDD_Mp9@2867_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2866 N_OUT9_Mp9@2866_d N_OUT8_Mp9@2866_g N_VDD_Mp9@2866_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2865 N_OUT9_Mn9@2865_d N_OUT8_Mn9@2865_g N_VSS_Mn9@2865_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2864 N_OUT9_Mn9@2864_d N_OUT8_Mn9@2864_g N_VSS_Mn9@2864_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2865 N_OUT9_Mp9@2865_d N_OUT8_Mp9@2865_g N_VDD_Mp9@2865_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2864 N_OUT9_Mp9@2864_d N_OUT8_Mp9@2864_g N_VDD_Mp9@2864_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2863 N_OUT9_Mn9@2863_d N_OUT8_Mn9@2863_g N_VSS_Mn9@2863_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2862 N_OUT9_Mn9@2862_d N_OUT8_Mn9@2862_g N_VSS_Mn9@2862_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2863 N_OUT9_Mp9@2863_d N_OUT8_Mp9@2863_g N_VDD_Mp9@2863_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2862 N_OUT9_Mp9@2862_d N_OUT8_Mp9@2862_g N_VDD_Mp9@2862_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2861 N_OUT9_Mn9@2861_d N_OUT8_Mn9@2861_g N_VSS_Mn9@2861_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2860 N_OUT9_Mn9@2860_d N_OUT8_Mn9@2860_g N_VSS_Mn9@2860_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2861 N_OUT9_Mp9@2861_d N_OUT8_Mp9@2861_g N_VDD_Mp9@2861_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2860 N_OUT9_Mp9@2860_d N_OUT8_Mp9@2860_g N_VDD_Mp9@2860_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2859 N_OUT9_Mn9@2859_d N_OUT8_Mn9@2859_g N_VSS_Mn9@2859_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2858 N_OUT9_Mn9@2858_d N_OUT8_Mn9@2858_g N_VSS_Mn9@2858_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2859 N_OUT9_Mp9@2859_d N_OUT8_Mp9@2859_g N_VDD_Mp9@2859_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2858 N_OUT9_Mp9@2858_d N_OUT8_Mp9@2858_g N_VDD_Mp9@2858_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2857 N_OUT9_Mn9@2857_d N_OUT8_Mn9@2857_g N_VSS_Mn9@2857_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2856 N_OUT9_Mn9@2856_d N_OUT8_Mn9@2856_g N_VSS_Mn9@2856_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2857 N_OUT9_Mp9@2857_d N_OUT8_Mp9@2857_g N_VDD_Mp9@2857_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2856 N_OUT9_Mp9@2856_d N_OUT8_Mp9@2856_g N_VDD_Mp9@2856_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2855 N_OUT9_Mn9@2855_d N_OUT8_Mn9@2855_g N_VSS_Mn9@2855_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2854 N_OUT9_Mn9@2854_d N_OUT8_Mn9@2854_g N_VSS_Mn9@2854_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2855 N_OUT9_Mp9@2855_d N_OUT8_Mp9@2855_g N_VDD_Mp9@2855_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2854 N_OUT9_Mp9@2854_d N_OUT8_Mp9@2854_g N_VDD_Mp9@2854_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2853 N_OUT9_Mn9@2853_d N_OUT8_Mn9@2853_g N_VSS_Mn9@2853_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2852 N_OUT9_Mn9@2852_d N_OUT8_Mn9@2852_g N_VSS_Mn9@2852_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2853 N_OUT9_Mp9@2853_d N_OUT8_Mp9@2853_g N_VDD_Mp9@2853_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2852 N_OUT9_Mp9@2852_d N_OUT8_Mp9@2852_g N_VDD_Mp9@2852_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2851 N_OUT9_Mn9@2851_d N_OUT8_Mn9@2851_g N_VSS_Mn9@2851_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2850 N_OUT9_Mn9@2850_d N_OUT8_Mn9@2850_g N_VSS_Mn9@2850_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2851 N_OUT9_Mp9@2851_d N_OUT8_Mp9@2851_g N_VDD_Mp9@2851_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2850 N_OUT9_Mp9@2850_d N_OUT8_Mp9@2850_g N_VDD_Mp9@2850_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2849 N_OUT9_Mn9@2849_d N_OUT8_Mn9@2849_g N_VSS_Mn9@2849_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2848 N_OUT9_Mn9@2848_d N_OUT8_Mn9@2848_g N_VSS_Mn9@2848_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2849 N_OUT9_Mp9@2849_d N_OUT8_Mp9@2849_g N_VDD_Mp9@2849_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2848 N_OUT9_Mp9@2848_d N_OUT8_Mp9@2848_g N_VDD_Mp9@2848_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2847 N_OUT9_Mn9@2847_d N_OUT8_Mn9@2847_g N_VSS_Mn9@2847_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2846 N_OUT9_Mn9@2846_d N_OUT8_Mn9@2846_g N_VSS_Mn9@2846_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2847 N_OUT9_Mp9@2847_d N_OUT8_Mp9@2847_g N_VDD_Mp9@2847_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2846 N_OUT9_Mp9@2846_d N_OUT8_Mp9@2846_g N_VDD_Mp9@2846_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2845 N_OUT9_Mn9@2845_d N_OUT8_Mn9@2845_g N_VSS_Mn9@2845_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2844 N_OUT9_Mn9@2844_d N_OUT8_Mn9@2844_g N_VSS_Mn9@2844_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2845 N_OUT9_Mp9@2845_d N_OUT8_Mp9@2845_g N_VDD_Mp9@2845_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2844 N_OUT9_Mp9@2844_d N_OUT8_Mp9@2844_g N_VDD_Mp9@2844_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2843 N_OUT9_Mn9@2843_d N_OUT8_Mn9@2843_g N_VSS_Mn9@2843_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2842 N_OUT9_Mn9@2842_d N_OUT8_Mn9@2842_g N_VSS_Mn9@2842_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2843 N_OUT9_Mp9@2843_d N_OUT8_Mp9@2843_g N_VDD_Mp9@2843_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2842 N_OUT9_Mp9@2842_d N_OUT8_Mp9@2842_g N_VDD_Mp9@2842_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2841 N_OUT9_Mn9@2841_d N_OUT8_Mn9@2841_g N_VSS_Mn9@2841_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2840 N_OUT9_Mn9@2840_d N_OUT8_Mn9@2840_g N_VSS_Mn9@2840_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2841 N_OUT9_Mp9@2841_d N_OUT8_Mp9@2841_g N_VDD_Mp9@2841_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2840 N_OUT9_Mp9@2840_d N_OUT8_Mp9@2840_g N_VDD_Mp9@2840_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2839 N_OUT9_Mn9@2839_d N_OUT8_Mn9@2839_g N_VSS_Mn9@2839_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2838 N_OUT9_Mn9@2838_d N_OUT8_Mn9@2838_g N_VSS_Mn9@2838_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2839 N_OUT9_Mp9@2839_d N_OUT8_Mp9@2839_g N_VDD_Mp9@2839_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2838 N_OUT9_Mp9@2838_d N_OUT8_Mp9@2838_g N_VDD_Mp9@2838_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2837 N_OUT9_Mn9@2837_d N_OUT8_Mn9@2837_g N_VSS_Mn9@2837_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2836 N_OUT9_Mn9@2836_d N_OUT8_Mn9@2836_g N_VSS_Mn9@2836_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2837 N_OUT9_Mp9@2837_d N_OUT8_Mp9@2837_g N_VDD_Mp9@2837_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2836 N_OUT9_Mp9@2836_d N_OUT8_Mp9@2836_g N_VDD_Mp9@2836_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2835 N_OUT9_Mn9@2835_d N_OUT8_Mn9@2835_g N_VSS_Mn9@2835_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2834 N_OUT9_Mn9@2834_d N_OUT8_Mn9@2834_g N_VSS_Mn9@2834_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2835 N_OUT9_Mp9@2835_d N_OUT8_Mp9@2835_g N_VDD_Mp9@2835_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2834 N_OUT9_Mp9@2834_d N_OUT8_Mp9@2834_g N_VDD_Mp9@2834_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2833 N_OUT9_Mn9@2833_d N_OUT8_Mn9@2833_g N_VSS_Mn9@2833_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2832 N_OUT9_Mn9@2832_d N_OUT8_Mn9@2832_g N_VSS_Mn9@2832_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2833 N_OUT9_Mp9@2833_d N_OUT8_Mp9@2833_g N_VDD_Mp9@2833_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2832 N_OUT9_Mp9@2832_d N_OUT8_Mp9@2832_g N_VDD_Mp9@2832_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2831 N_OUT9_Mn9@2831_d N_OUT8_Mn9@2831_g N_VSS_Mn9@2831_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2830 N_OUT9_Mn9@2830_d N_OUT8_Mn9@2830_g N_VSS_Mn9@2830_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2831 N_OUT9_Mp9@2831_d N_OUT8_Mp9@2831_g N_VDD_Mp9@2831_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2830 N_OUT9_Mp9@2830_d N_OUT8_Mp9@2830_g N_VDD_Mp9@2830_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2829 N_OUT9_Mn9@2829_d N_OUT8_Mn9@2829_g N_VSS_Mn9@2829_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2828 N_OUT9_Mn9@2828_d N_OUT8_Mn9@2828_g N_VSS_Mn9@2828_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2829 N_OUT9_Mp9@2829_d N_OUT8_Mp9@2829_g N_VDD_Mp9@2829_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2828 N_OUT9_Mp9@2828_d N_OUT8_Mp9@2828_g N_VDD_Mp9@2828_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2827 N_OUT9_Mn9@2827_d N_OUT8_Mn9@2827_g N_VSS_Mn9@2827_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2826 N_OUT9_Mn9@2826_d N_OUT8_Mn9@2826_g N_VSS_Mn9@2826_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2827 N_OUT9_Mp9@2827_d N_OUT8_Mp9@2827_g N_VDD_Mp9@2827_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2826 N_OUT9_Mp9@2826_d N_OUT8_Mp9@2826_g N_VDD_Mp9@2826_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2825 N_OUT9_Mn9@2825_d N_OUT8_Mn9@2825_g N_VSS_Mn9@2825_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2824 N_OUT9_Mn9@2824_d N_OUT8_Mn9@2824_g N_VSS_Mn9@2824_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2825 N_OUT9_Mp9@2825_d N_OUT8_Mp9@2825_g N_VDD_Mp9@2825_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2824 N_OUT9_Mp9@2824_d N_OUT8_Mp9@2824_g N_VDD_Mp9@2824_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2823 N_OUT9_Mn9@2823_d N_OUT8_Mn9@2823_g N_VSS_Mn9@2823_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2822 N_OUT9_Mn9@2822_d N_OUT8_Mn9@2822_g N_VSS_Mn9@2822_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2823 N_OUT9_Mp9@2823_d N_OUT8_Mp9@2823_g N_VDD_Mp9@2823_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2822 N_OUT9_Mp9@2822_d N_OUT8_Mp9@2822_g N_VDD_Mp9@2822_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2821 N_OUT9_Mn9@2821_d N_OUT8_Mn9@2821_g N_VSS_Mn9@2821_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2820 N_OUT9_Mn9@2820_d N_OUT8_Mn9@2820_g N_VSS_Mn9@2820_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2821 N_OUT9_Mp9@2821_d N_OUT8_Mp9@2821_g N_VDD_Mp9@2821_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2820 N_OUT9_Mp9@2820_d N_OUT8_Mp9@2820_g N_VDD_Mp9@2820_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2819 N_OUT9_Mn9@2819_d N_OUT8_Mn9@2819_g N_VSS_Mn9@2819_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2818 N_OUT9_Mn9@2818_d N_OUT8_Mn9@2818_g N_VSS_Mn9@2818_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2819 N_OUT9_Mp9@2819_d N_OUT8_Mp9@2819_g N_VDD_Mp9@2819_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2818 N_OUT9_Mp9@2818_d N_OUT8_Mp9@2818_g N_VDD_Mp9@2818_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2817 N_OUT9_Mn9@2817_d N_OUT8_Mn9@2817_g N_VSS_Mn9@2817_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2816 N_OUT9_Mn9@2816_d N_OUT8_Mn9@2816_g N_VSS_Mn9@2816_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2817 N_OUT9_Mp9@2817_d N_OUT8_Mp9@2817_g N_VDD_Mp9@2817_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2816 N_OUT9_Mp9@2816_d N_OUT8_Mp9@2816_g N_VDD_Mp9@2816_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2815 N_OUT9_Mn9@2815_d N_OUT8_Mn9@2815_g N_VSS_Mn9@2815_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2814 N_OUT9_Mn9@2814_d N_OUT8_Mn9@2814_g N_VSS_Mn9@2814_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2815 N_OUT9_Mp9@2815_d N_OUT8_Mp9@2815_g N_VDD_Mp9@2815_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2814 N_OUT9_Mp9@2814_d N_OUT8_Mp9@2814_g N_VDD_Mp9@2814_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2813 N_OUT9_Mn9@2813_d N_OUT8_Mn9@2813_g N_VSS_Mn9@2813_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2812 N_OUT9_Mn9@2812_d N_OUT8_Mn9@2812_g N_VSS_Mn9@2812_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2813 N_OUT9_Mp9@2813_d N_OUT8_Mp9@2813_g N_VDD_Mp9@2813_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2812 N_OUT9_Mp9@2812_d N_OUT8_Mp9@2812_g N_VDD_Mp9@2812_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2811 N_OUT9_Mn9@2811_d N_OUT8_Mn9@2811_g N_VSS_Mn9@2811_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2810 N_OUT9_Mn9@2810_d N_OUT8_Mn9@2810_g N_VSS_Mn9@2810_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2811 N_OUT9_Mp9@2811_d N_OUT8_Mp9@2811_g N_VDD_Mp9@2811_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2810 N_OUT9_Mp9@2810_d N_OUT8_Mp9@2810_g N_VDD_Mp9@2810_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2809 N_OUT9_Mn9@2809_d N_OUT8_Mn9@2809_g N_VSS_Mn9@2809_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2808 N_OUT9_Mn9@2808_d N_OUT8_Mn9@2808_g N_VSS_Mn9@2808_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2809 N_OUT9_Mp9@2809_d N_OUT8_Mp9@2809_g N_VDD_Mp9@2809_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2808 N_OUT9_Mp9@2808_d N_OUT8_Mp9@2808_g N_VDD_Mp9@2808_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2807 N_OUT9_Mn9@2807_d N_OUT8_Mn9@2807_g N_VSS_Mn9@2807_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2806 N_OUT9_Mn9@2806_d N_OUT8_Mn9@2806_g N_VSS_Mn9@2806_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2807 N_OUT9_Mp9@2807_d N_OUT8_Mp9@2807_g N_VDD_Mp9@2807_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2806 N_OUT9_Mp9@2806_d N_OUT8_Mp9@2806_g N_VDD_Mp9@2806_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2805 N_OUT9_Mn9@2805_d N_OUT8_Mn9@2805_g N_VSS_Mn9@2805_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2804 N_OUT9_Mn9@2804_d N_OUT8_Mn9@2804_g N_VSS_Mn9@2804_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2805 N_OUT9_Mp9@2805_d N_OUT8_Mp9@2805_g N_VDD_Mp9@2805_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2804 N_OUT9_Mp9@2804_d N_OUT8_Mp9@2804_g N_VDD_Mp9@2804_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2803 N_OUT9_Mn9@2803_d N_OUT8_Mn9@2803_g N_VSS_Mn9@2803_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2802 N_OUT9_Mn9@2802_d N_OUT8_Mn9@2802_g N_VSS_Mn9@2802_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2803 N_OUT9_Mp9@2803_d N_OUT8_Mp9@2803_g N_VDD_Mp9@2803_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2802 N_OUT9_Mp9@2802_d N_OUT8_Mp9@2802_g N_VDD_Mp9@2802_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2801 N_OUT9_Mn9@2801_d N_OUT8_Mn9@2801_g N_VSS_Mn9@2801_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2800 N_OUT9_Mn9@2800_d N_OUT8_Mn9@2800_g N_VSS_Mn9@2800_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2801 N_OUT9_Mp9@2801_d N_OUT8_Mp9@2801_g N_VDD_Mp9@2801_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2800 N_OUT9_Mp9@2800_d N_OUT8_Mp9@2800_g N_VDD_Mp9@2800_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2799 N_OUT9_Mn9@2799_d N_OUT8_Mn9@2799_g N_VSS_Mn9@2799_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2798 N_OUT9_Mn9@2798_d N_OUT8_Mn9@2798_g N_VSS_Mn9@2798_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2799 N_OUT9_Mp9@2799_d N_OUT8_Mp9@2799_g N_VDD_Mp9@2799_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2798 N_OUT9_Mp9@2798_d N_OUT8_Mp9@2798_g N_VDD_Mp9@2798_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2797 N_OUT9_Mn9@2797_d N_OUT8_Mn9@2797_g N_VSS_Mn9@2797_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2796 N_OUT9_Mn9@2796_d N_OUT8_Mn9@2796_g N_VSS_Mn9@2796_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2797 N_OUT9_Mp9@2797_d N_OUT8_Mp9@2797_g N_VDD_Mp9@2797_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2796 N_OUT9_Mp9@2796_d N_OUT8_Mp9@2796_g N_VDD_Mp9@2796_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2795 N_OUT9_Mn9@2795_d N_OUT8_Mn9@2795_g N_VSS_Mn9@2795_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2794 N_OUT9_Mn9@2794_d N_OUT8_Mn9@2794_g N_VSS_Mn9@2794_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2795 N_OUT9_Mp9@2795_d N_OUT8_Mp9@2795_g N_VDD_Mp9@2795_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2794 N_OUT9_Mp9@2794_d N_OUT8_Mp9@2794_g N_VDD_Mp9@2794_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2793 N_OUT9_Mn9@2793_d N_OUT8_Mn9@2793_g N_VSS_Mn9@2793_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2792 N_OUT9_Mn9@2792_d N_OUT8_Mn9@2792_g N_VSS_Mn9@2792_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2793 N_OUT9_Mp9@2793_d N_OUT8_Mp9@2793_g N_VDD_Mp9@2793_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2792 N_OUT9_Mp9@2792_d N_OUT8_Mp9@2792_g N_VDD_Mp9@2792_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2791 N_OUT9_Mn9@2791_d N_OUT8_Mn9@2791_g N_VSS_Mn9@2791_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2790 N_OUT9_Mn9@2790_d N_OUT8_Mn9@2790_g N_VSS_Mn9@2790_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2791 N_OUT9_Mp9@2791_d N_OUT8_Mp9@2791_g N_VDD_Mp9@2791_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2790 N_OUT9_Mp9@2790_d N_OUT8_Mp9@2790_g N_VDD_Mp9@2790_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2789 N_OUT9_Mn9@2789_d N_OUT8_Mn9@2789_g N_VSS_Mn9@2789_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2788 N_OUT9_Mn9@2788_d N_OUT8_Mn9@2788_g N_VSS_Mn9@2788_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2789 N_OUT9_Mp9@2789_d N_OUT8_Mp9@2789_g N_VDD_Mp9@2789_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2788 N_OUT9_Mp9@2788_d N_OUT8_Mp9@2788_g N_VDD_Mp9@2788_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2787 N_OUT9_Mn9@2787_d N_OUT8_Mn9@2787_g N_VSS_Mn9@2787_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2786 N_OUT9_Mn9@2786_d N_OUT8_Mn9@2786_g N_VSS_Mn9@2786_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2787 N_OUT9_Mp9@2787_d N_OUT8_Mp9@2787_g N_VDD_Mp9@2787_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2786 N_OUT9_Mp9@2786_d N_OUT8_Mp9@2786_g N_VDD_Mp9@2786_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2785 N_OUT9_Mn9@2785_d N_OUT8_Mn9@2785_g N_VSS_Mn9@2785_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2784 N_OUT9_Mn9@2784_d N_OUT8_Mn9@2784_g N_VSS_Mn9@2784_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2785 N_OUT9_Mp9@2785_d N_OUT8_Mp9@2785_g N_VDD_Mp9@2785_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2784 N_OUT9_Mp9@2784_d N_OUT8_Mp9@2784_g N_VDD_Mp9@2784_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2783 N_OUT9_Mn9@2783_d N_OUT8_Mn9@2783_g N_VSS_Mn9@2783_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2782 N_OUT9_Mn9@2782_d N_OUT8_Mn9@2782_g N_VSS_Mn9@2782_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2783 N_OUT9_Mp9@2783_d N_OUT8_Mp9@2783_g N_VDD_Mp9@2783_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2782 N_OUT9_Mp9@2782_d N_OUT8_Mp9@2782_g N_VDD_Mp9@2782_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2781 N_OUT9_Mn9@2781_d N_OUT8_Mn9@2781_g N_VSS_Mn9@2781_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2780 N_OUT9_Mn9@2780_d N_OUT8_Mn9@2780_g N_VSS_Mn9@2780_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2781 N_OUT9_Mp9@2781_d N_OUT8_Mp9@2781_g N_VDD_Mp9@2781_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2780 N_OUT9_Mp9@2780_d N_OUT8_Mp9@2780_g N_VDD_Mp9@2780_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2779 N_OUT9_Mn9@2779_d N_OUT8_Mn9@2779_g N_VSS_Mn9@2779_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2778 N_OUT9_Mn9@2778_d N_OUT8_Mn9@2778_g N_VSS_Mn9@2778_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2779 N_OUT9_Mp9@2779_d N_OUT8_Mp9@2779_g N_VDD_Mp9@2779_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2778 N_OUT9_Mp9@2778_d N_OUT8_Mp9@2778_g N_VDD_Mp9@2778_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2777 N_OUT9_Mn9@2777_d N_OUT8_Mn9@2777_g N_VSS_Mn9@2777_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2776 N_OUT9_Mn9@2776_d N_OUT8_Mn9@2776_g N_VSS_Mn9@2776_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2777 N_OUT9_Mp9@2777_d N_OUT8_Mp9@2777_g N_VDD_Mp9@2777_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2776 N_OUT9_Mp9@2776_d N_OUT8_Mp9@2776_g N_VDD_Mp9@2776_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2775 N_OUT9_Mn9@2775_d N_OUT8_Mn9@2775_g N_VSS_Mn9@2775_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2774 N_OUT9_Mn9@2774_d N_OUT8_Mn9@2774_g N_VSS_Mn9@2774_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2775 N_OUT9_Mp9@2775_d N_OUT8_Mp9@2775_g N_VDD_Mp9@2775_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2774 N_OUT9_Mp9@2774_d N_OUT8_Mp9@2774_g N_VDD_Mp9@2774_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2773 N_OUT9_Mn9@2773_d N_OUT8_Mn9@2773_g N_VSS_Mn9@2773_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2772 N_OUT9_Mn9@2772_d N_OUT8_Mn9@2772_g N_VSS_Mn9@2772_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2773 N_OUT9_Mp9@2773_d N_OUT8_Mp9@2773_g N_VDD_Mp9@2773_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2772 N_OUT9_Mp9@2772_d N_OUT8_Mp9@2772_g N_VDD_Mp9@2772_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2771 N_OUT9_Mn9@2771_d N_OUT8_Mn9@2771_g N_VSS_Mn9@2771_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2770 N_OUT9_Mn9@2770_d N_OUT8_Mn9@2770_g N_VSS_Mn9@2770_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2771 N_OUT9_Mp9@2771_d N_OUT8_Mp9@2771_g N_VDD_Mp9@2771_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2770 N_OUT9_Mp9@2770_d N_OUT8_Mp9@2770_g N_VDD_Mp9@2770_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2769 N_OUT9_Mn9@2769_d N_OUT8_Mn9@2769_g N_VSS_Mn9@2769_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2768 N_OUT9_Mn9@2768_d N_OUT8_Mn9@2768_g N_VSS_Mn9@2768_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2769 N_OUT9_Mp9@2769_d N_OUT8_Mp9@2769_g N_VDD_Mp9@2769_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2768 N_OUT9_Mp9@2768_d N_OUT8_Mp9@2768_g N_VDD_Mp9@2768_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2767 N_OUT9_Mn9@2767_d N_OUT8_Mn9@2767_g N_VSS_Mn9@2767_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2766 N_OUT9_Mn9@2766_d N_OUT8_Mn9@2766_g N_VSS_Mn9@2766_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2767 N_OUT9_Mp9@2767_d N_OUT8_Mp9@2767_g N_VDD_Mp9@2767_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2766 N_OUT9_Mp9@2766_d N_OUT8_Mp9@2766_g N_VDD_Mp9@2766_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2765 N_OUT9_Mn9@2765_d N_OUT8_Mn9@2765_g N_VSS_Mn9@2765_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2764 N_OUT9_Mn9@2764_d N_OUT8_Mn9@2764_g N_VSS_Mn9@2764_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2765 N_OUT9_Mp9@2765_d N_OUT8_Mp9@2765_g N_VDD_Mp9@2765_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2764 N_OUT9_Mp9@2764_d N_OUT8_Mp9@2764_g N_VDD_Mp9@2764_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2763 N_OUT9_Mn9@2763_d N_OUT8_Mn9@2763_g N_VSS_Mn9@2763_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2762 N_OUT9_Mn9@2762_d N_OUT8_Mn9@2762_g N_VSS_Mn9@2762_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2763 N_OUT9_Mp9@2763_d N_OUT8_Mp9@2763_g N_VDD_Mp9@2763_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2762 N_OUT9_Mp9@2762_d N_OUT8_Mp9@2762_g N_VDD_Mp9@2762_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2761 N_OUT9_Mn9@2761_d N_OUT8_Mn9@2761_g N_VSS_Mn9@2761_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2760 N_OUT9_Mn9@2760_d N_OUT8_Mn9@2760_g N_VSS_Mn9@2760_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2761 N_OUT9_Mp9@2761_d N_OUT8_Mp9@2761_g N_VDD_Mp9@2761_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2760 N_OUT9_Mp9@2760_d N_OUT8_Mp9@2760_g N_VDD_Mp9@2760_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2759 N_OUT9_Mn9@2759_d N_OUT8_Mn9@2759_g N_VSS_Mn9@2759_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2758 N_OUT9_Mn9@2758_d N_OUT8_Mn9@2758_g N_VSS_Mn9@2758_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2759 N_OUT9_Mp9@2759_d N_OUT8_Mp9@2759_g N_VDD_Mp9@2759_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2758 N_OUT9_Mp9@2758_d N_OUT8_Mp9@2758_g N_VDD_Mp9@2758_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2757 N_OUT9_Mn9@2757_d N_OUT8_Mn9@2757_g N_VSS_Mn9@2757_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2756 N_OUT9_Mn9@2756_d N_OUT8_Mn9@2756_g N_VSS_Mn9@2756_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2757 N_OUT9_Mp9@2757_d N_OUT8_Mp9@2757_g N_VDD_Mp9@2757_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2756 N_OUT9_Mp9@2756_d N_OUT8_Mp9@2756_g N_VDD_Mp9@2756_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2755 N_OUT9_Mn9@2755_d N_OUT8_Mn9@2755_g N_VSS_Mn9@2755_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2754 N_OUT9_Mn9@2754_d N_OUT8_Mn9@2754_g N_VSS_Mn9@2754_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2755 N_OUT9_Mp9@2755_d N_OUT8_Mp9@2755_g N_VDD_Mp9@2755_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2754 N_OUT9_Mp9@2754_d N_OUT8_Mp9@2754_g N_VDD_Mp9@2754_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2753 N_OUT9_Mn9@2753_d N_OUT8_Mn9@2753_g N_VSS_Mn9@2753_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2752 N_OUT9_Mn9@2752_d N_OUT8_Mn9@2752_g N_VSS_Mn9@2752_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2753 N_OUT9_Mp9@2753_d N_OUT8_Mp9@2753_g N_VDD_Mp9@2753_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2752 N_OUT9_Mp9@2752_d N_OUT8_Mp9@2752_g N_VDD_Mp9@2752_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2751 N_OUT9_Mn9@2751_d N_OUT8_Mn9@2751_g N_VSS_Mn9@2751_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2750 N_OUT9_Mn9@2750_d N_OUT8_Mn9@2750_g N_VSS_Mn9@2750_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2751 N_OUT9_Mp9@2751_d N_OUT8_Mp9@2751_g N_VDD_Mp9@2751_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2750 N_OUT9_Mp9@2750_d N_OUT8_Mp9@2750_g N_VDD_Mp9@2750_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2749 N_OUT9_Mn9@2749_d N_OUT8_Mn9@2749_g N_VSS_Mn9@2749_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2748 N_OUT9_Mn9@2748_d N_OUT8_Mn9@2748_g N_VSS_Mn9@2748_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2749 N_OUT9_Mp9@2749_d N_OUT8_Mp9@2749_g N_VDD_Mp9@2749_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2748 N_OUT9_Mp9@2748_d N_OUT8_Mp9@2748_g N_VDD_Mp9@2748_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2747 N_OUT9_Mn9@2747_d N_OUT8_Mn9@2747_g N_VSS_Mn9@2747_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2746 N_OUT9_Mn9@2746_d N_OUT8_Mn9@2746_g N_VSS_Mn9@2746_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2747 N_OUT9_Mp9@2747_d N_OUT8_Mp9@2747_g N_VDD_Mp9@2747_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2746 N_OUT9_Mp9@2746_d N_OUT8_Mp9@2746_g N_VDD_Mp9@2746_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2745 N_OUT9_Mn9@2745_d N_OUT8_Mn9@2745_g N_VSS_Mn9@2745_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2744 N_OUT9_Mn9@2744_d N_OUT8_Mn9@2744_g N_VSS_Mn9@2744_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2745 N_OUT9_Mp9@2745_d N_OUT8_Mp9@2745_g N_VDD_Mp9@2745_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2744 N_OUT9_Mp9@2744_d N_OUT8_Mp9@2744_g N_VDD_Mp9@2744_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2743 N_OUT9_Mn9@2743_d N_OUT8_Mn9@2743_g N_VSS_Mn9@2743_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2742 N_OUT9_Mn9@2742_d N_OUT8_Mn9@2742_g N_VSS_Mn9@2742_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2743 N_OUT9_Mp9@2743_d N_OUT8_Mp9@2743_g N_VDD_Mp9@2743_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2742 N_OUT9_Mp9@2742_d N_OUT8_Mp9@2742_g N_VDD_Mp9@2742_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2741 N_OUT9_Mn9@2741_d N_OUT8_Mn9@2741_g N_VSS_Mn9@2741_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2740 N_OUT9_Mn9@2740_d N_OUT8_Mn9@2740_g N_VSS_Mn9@2740_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2741 N_OUT9_Mp9@2741_d N_OUT8_Mp9@2741_g N_VDD_Mp9@2741_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2740 N_OUT9_Mp9@2740_d N_OUT8_Mp9@2740_g N_VDD_Mp9@2740_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2739 N_OUT9_Mn9@2739_d N_OUT8_Mn9@2739_g N_VSS_Mn9@2739_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2738 N_OUT9_Mn9@2738_d N_OUT8_Mn9@2738_g N_VSS_Mn9@2738_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2739 N_OUT9_Mp9@2739_d N_OUT8_Mp9@2739_g N_VDD_Mp9@2739_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2738 N_OUT9_Mp9@2738_d N_OUT8_Mp9@2738_g N_VDD_Mp9@2738_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2737 N_OUT9_Mn9@2737_d N_OUT8_Mn9@2737_g N_VSS_Mn9@2737_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2736 N_OUT9_Mn9@2736_d N_OUT8_Mn9@2736_g N_VSS_Mn9@2736_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2737 N_OUT9_Mp9@2737_d N_OUT8_Mp9@2737_g N_VDD_Mp9@2737_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2736 N_OUT9_Mp9@2736_d N_OUT8_Mp9@2736_g N_VDD_Mp9@2736_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2735 N_OUT9_Mn9@2735_d N_OUT8_Mn9@2735_g N_VSS_Mn9@2735_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2734 N_OUT9_Mn9@2734_d N_OUT8_Mn9@2734_g N_VSS_Mn9@2734_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2735 N_OUT9_Mp9@2735_d N_OUT8_Mp9@2735_g N_VDD_Mp9@2735_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2734 N_OUT9_Mp9@2734_d N_OUT8_Mp9@2734_g N_VDD_Mp9@2734_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2733 N_OUT9_Mn9@2733_d N_OUT8_Mn9@2733_g N_VSS_Mn9@2733_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2732 N_OUT9_Mn9@2732_d N_OUT8_Mn9@2732_g N_VSS_Mn9@2732_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2733 N_OUT9_Mp9@2733_d N_OUT8_Mp9@2733_g N_VDD_Mp9@2733_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2732 N_OUT9_Mp9@2732_d N_OUT8_Mp9@2732_g N_VDD_Mp9@2732_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2731 N_OUT9_Mn9@2731_d N_OUT8_Mn9@2731_g N_VSS_Mn9@2731_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2730 N_OUT9_Mn9@2730_d N_OUT8_Mn9@2730_g N_VSS_Mn9@2730_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2731 N_OUT9_Mp9@2731_d N_OUT8_Mp9@2731_g N_VDD_Mp9@2731_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2730 N_OUT9_Mp9@2730_d N_OUT8_Mp9@2730_g N_VDD_Mp9@2730_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2729 N_OUT9_Mn9@2729_d N_OUT8_Mn9@2729_g N_VSS_Mn9@2729_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2728 N_OUT9_Mn9@2728_d N_OUT8_Mn9@2728_g N_VSS_Mn9@2728_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2729 N_OUT9_Mp9@2729_d N_OUT8_Mp9@2729_g N_VDD_Mp9@2729_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2728 N_OUT9_Mp9@2728_d N_OUT8_Mp9@2728_g N_VDD_Mp9@2728_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2727 N_OUT9_Mn9@2727_d N_OUT8_Mn9@2727_g N_VSS_Mn9@2727_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2726 N_OUT9_Mn9@2726_d N_OUT8_Mn9@2726_g N_VSS_Mn9@2726_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2727 N_OUT9_Mp9@2727_d N_OUT8_Mp9@2727_g N_VDD_Mp9@2727_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2726 N_OUT9_Mp9@2726_d N_OUT8_Mp9@2726_g N_VDD_Mp9@2726_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2725 N_OUT9_Mn9@2725_d N_OUT8_Mn9@2725_g N_VSS_Mn9@2725_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2724 N_OUT9_Mn9@2724_d N_OUT8_Mn9@2724_g N_VSS_Mn9@2724_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2725 N_OUT9_Mp9@2725_d N_OUT8_Mp9@2725_g N_VDD_Mp9@2725_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2724 N_OUT9_Mp9@2724_d N_OUT8_Mp9@2724_g N_VDD_Mp9@2724_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2723 N_OUT9_Mn9@2723_d N_OUT8_Mn9@2723_g N_VSS_Mn9@2723_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2722 N_OUT9_Mn9@2722_d N_OUT8_Mn9@2722_g N_VSS_Mn9@2722_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2723 N_OUT9_Mp9@2723_d N_OUT8_Mp9@2723_g N_VDD_Mp9@2723_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2722 N_OUT9_Mp9@2722_d N_OUT8_Mp9@2722_g N_VDD_Mp9@2722_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2721 N_OUT9_Mn9@2721_d N_OUT8_Mn9@2721_g N_VSS_Mn9@2721_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2720 N_OUT9_Mn9@2720_d N_OUT8_Mn9@2720_g N_VSS_Mn9@2720_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2721 N_OUT9_Mp9@2721_d N_OUT8_Mp9@2721_g N_VDD_Mp9@2721_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2720 N_OUT9_Mp9@2720_d N_OUT8_Mp9@2720_g N_VDD_Mp9@2720_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2719 N_OUT9_Mn9@2719_d N_OUT8_Mn9@2719_g N_VSS_Mn9@2719_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2718 N_OUT9_Mn9@2718_d N_OUT8_Mn9@2718_g N_VSS_Mn9@2718_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2719 N_OUT9_Mp9@2719_d N_OUT8_Mp9@2719_g N_VDD_Mp9@2719_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2718 N_OUT9_Mp9@2718_d N_OUT8_Mp9@2718_g N_VDD_Mp9@2718_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2717 N_OUT9_Mn9@2717_d N_OUT8_Mn9@2717_g N_VSS_Mn9@2717_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2716 N_OUT9_Mn9@2716_d N_OUT8_Mn9@2716_g N_VSS_Mn9@2716_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2717 N_OUT9_Mp9@2717_d N_OUT8_Mp9@2717_g N_VDD_Mp9@2717_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2716 N_OUT9_Mp9@2716_d N_OUT8_Mp9@2716_g N_VDD_Mp9@2716_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2715 N_OUT9_Mn9@2715_d N_OUT8_Mn9@2715_g N_VSS_Mn9@2715_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2714 N_OUT9_Mn9@2714_d N_OUT8_Mn9@2714_g N_VSS_Mn9@2714_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2715 N_OUT9_Mp9@2715_d N_OUT8_Mp9@2715_g N_VDD_Mp9@2715_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2714 N_OUT9_Mp9@2714_d N_OUT8_Mp9@2714_g N_VDD_Mp9@2714_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2713 N_OUT9_Mn9@2713_d N_OUT8_Mn9@2713_g N_VSS_Mn9@2713_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2712 N_OUT9_Mn9@2712_d N_OUT8_Mn9@2712_g N_VSS_Mn9@2712_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2713 N_OUT9_Mp9@2713_d N_OUT8_Mp9@2713_g N_VDD_Mp9@2713_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2712 N_OUT9_Mp9@2712_d N_OUT8_Mp9@2712_g N_VDD_Mp9@2712_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2711 N_OUT9_Mn9@2711_d N_OUT8_Mn9@2711_g N_VSS_Mn9@2711_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2710 N_OUT9_Mn9@2710_d N_OUT8_Mn9@2710_g N_VSS_Mn9@2710_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2711 N_OUT9_Mp9@2711_d N_OUT8_Mp9@2711_g N_VDD_Mp9@2711_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2710 N_OUT9_Mp9@2710_d N_OUT8_Mp9@2710_g N_VDD_Mp9@2710_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2709 N_OUT9_Mn9@2709_d N_OUT8_Mn9@2709_g N_VSS_Mn9@2709_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2708 N_OUT9_Mn9@2708_d N_OUT8_Mn9@2708_g N_VSS_Mn9@2708_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2709 N_OUT9_Mp9@2709_d N_OUT8_Mp9@2709_g N_VDD_Mp9@2709_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2708 N_OUT9_Mp9@2708_d N_OUT8_Mp9@2708_g N_VDD_Mp9@2708_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2707 N_OUT9_Mn9@2707_d N_OUT8_Mn9@2707_g N_VSS_Mn9@2707_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2706 N_OUT9_Mn9@2706_d N_OUT8_Mn9@2706_g N_VSS_Mn9@2706_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2707 N_OUT9_Mp9@2707_d N_OUT8_Mp9@2707_g N_VDD_Mp9@2707_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2706 N_OUT9_Mp9@2706_d N_OUT8_Mp9@2706_g N_VDD_Mp9@2706_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2705 N_OUT9_Mn9@2705_d N_OUT8_Mn9@2705_g N_VSS_Mn9@2705_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2704 N_OUT9_Mn9@2704_d N_OUT8_Mn9@2704_g N_VSS_Mn9@2704_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2705 N_OUT9_Mp9@2705_d N_OUT8_Mp9@2705_g N_VDD_Mp9@2705_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2704 N_OUT9_Mp9@2704_d N_OUT8_Mp9@2704_g N_VDD_Mp9@2704_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2703 N_OUT9_Mn9@2703_d N_OUT8_Mn9@2703_g N_VSS_Mn9@2703_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2702 N_OUT9_Mn9@2702_d N_OUT8_Mn9@2702_g N_VSS_Mn9@2702_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2703 N_OUT9_Mp9@2703_d N_OUT8_Mp9@2703_g N_VDD_Mp9@2703_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2702 N_OUT9_Mp9@2702_d N_OUT8_Mp9@2702_g N_VDD_Mp9@2702_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2701 N_OUT9_Mn9@2701_d N_OUT8_Mn9@2701_g N_VSS_Mn9@2701_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2700 N_OUT9_Mn9@2700_d N_OUT8_Mn9@2700_g N_VSS_Mn9@2700_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2701 N_OUT9_Mp9@2701_d N_OUT8_Mp9@2701_g N_VDD_Mp9@2701_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2700 N_OUT9_Mp9@2700_d N_OUT8_Mp9@2700_g N_VDD_Mp9@2700_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2699 N_OUT9_Mn9@2699_d N_OUT8_Mn9@2699_g N_VSS_Mn9@2699_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2698 N_OUT9_Mn9@2698_d N_OUT8_Mn9@2698_g N_VSS_Mn9@2698_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2699 N_OUT9_Mp9@2699_d N_OUT8_Mp9@2699_g N_VDD_Mp9@2699_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2698 N_OUT9_Mp9@2698_d N_OUT8_Mp9@2698_g N_VDD_Mp9@2698_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2697 N_OUT9_Mn9@2697_d N_OUT8_Mn9@2697_g N_VSS_Mn9@2697_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2696 N_OUT9_Mn9@2696_d N_OUT8_Mn9@2696_g N_VSS_Mn9@2696_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2697 N_OUT9_Mp9@2697_d N_OUT8_Mp9@2697_g N_VDD_Mp9@2697_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2696 N_OUT9_Mp9@2696_d N_OUT8_Mp9@2696_g N_VDD_Mp9@2696_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2695 N_OUT9_Mn9@2695_d N_OUT8_Mn9@2695_g N_VSS_Mn9@2695_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2694 N_OUT9_Mn9@2694_d N_OUT8_Mn9@2694_g N_VSS_Mn9@2694_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2695 N_OUT9_Mp9@2695_d N_OUT8_Mp9@2695_g N_VDD_Mp9@2695_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2694 N_OUT9_Mp9@2694_d N_OUT8_Mp9@2694_g N_VDD_Mp9@2694_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2693 N_OUT9_Mn9@2693_d N_OUT8_Mn9@2693_g N_VSS_Mn9@2693_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2692 N_OUT9_Mn9@2692_d N_OUT8_Mn9@2692_g N_VSS_Mn9@2692_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2693 N_OUT9_Mp9@2693_d N_OUT8_Mp9@2693_g N_VDD_Mp9@2693_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2692 N_OUT9_Mp9@2692_d N_OUT8_Mp9@2692_g N_VDD_Mp9@2692_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2691 N_OUT9_Mn9@2691_d N_OUT8_Mn9@2691_g N_VSS_Mn9@2691_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2690 N_OUT9_Mn9@2690_d N_OUT8_Mn9@2690_g N_VSS_Mn9@2690_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2691 N_OUT9_Mp9@2691_d N_OUT8_Mp9@2691_g N_VDD_Mp9@2691_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2690 N_OUT9_Mp9@2690_d N_OUT8_Mp9@2690_g N_VDD_Mp9@2690_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2689 N_OUT9_Mn9@2689_d N_OUT8_Mn9@2689_g N_VSS_Mn9@2689_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2688 N_OUT9_Mn9@2688_d N_OUT8_Mn9@2688_g N_VSS_Mn9@2688_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2689 N_OUT9_Mp9@2689_d N_OUT8_Mp9@2689_g N_VDD_Mp9@2689_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2688 N_OUT9_Mp9@2688_d N_OUT8_Mp9@2688_g N_VDD_Mp9@2688_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2687 N_OUT9_Mn9@2687_d N_OUT8_Mn9@2687_g N_VSS_Mn9@2687_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2686 N_OUT9_Mn9@2686_d N_OUT8_Mn9@2686_g N_VSS_Mn9@2686_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2687 N_OUT9_Mp9@2687_d N_OUT8_Mp9@2687_g N_VDD_Mp9@2687_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2686 N_OUT9_Mp9@2686_d N_OUT8_Mp9@2686_g N_VDD_Mp9@2686_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2685 N_OUT9_Mn9@2685_d N_OUT8_Mn9@2685_g N_VSS_Mn9@2685_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2684 N_OUT9_Mn9@2684_d N_OUT8_Mn9@2684_g N_VSS_Mn9@2684_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2685 N_OUT9_Mp9@2685_d N_OUT8_Mp9@2685_g N_VDD_Mp9@2685_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2684 N_OUT9_Mp9@2684_d N_OUT8_Mp9@2684_g N_VDD_Mp9@2684_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2683 N_OUT9_Mn9@2683_d N_OUT8_Mn9@2683_g N_VSS_Mn9@2683_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2682 N_OUT9_Mn9@2682_d N_OUT8_Mn9@2682_g N_VSS_Mn9@2682_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2683 N_OUT9_Mp9@2683_d N_OUT8_Mp9@2683_g N_VDD_Mp9@2683_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2682 N_OUT9_Mp9@2682_d N_OUT8_Mp9@2682_g N_VDD_Mp9@2682_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2681 N_OUT9_Mn9@2681_d N_OUT8_Mn9@2681_g N_VSS_Mn9@2681_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2680 N_OUT9_Mn9@2680_d N_OUT8_Mn9@2680_g N_VSS_Mn9@2680_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2681 N_OUT9_Mp9@2681_d N_OUT8_Mp9@2681_g N_VDD_Mp9@2681_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2680 N_OUT9_Mp9@2680_d N_OUT8_Mp9@2680_g N_VDD_Mp9@2680_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2679 N_OUT9_Mn9@2679_d N_OUT8_Mn9@2679_g N_VSS_Mn9@2679_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2678 N_OUT9_Mn9@2678_d N_OUT8_Mn9@2678_g N_VSS_Mn9@2678_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2679 N_OUT9_Mp9@2679_d N_OUT8_Mp9@2679_g N_VDD_Mp9@2679_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2678 N_OUT9_Mp9@2678_d N_OUT8_Mp9@2678_g N_VDD_Mp9@2678_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2677 N_OUT9_Mn9@2677_d N_OUT8_Mn9@2677_g N_VSS_Mn9@2677_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2676 N_OUT9_Mn9@2676_d N_OUT8_Mn9@2676_g N_VSS_Mn9@2676_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2677 N_OUT9_Mp9@2677_d N_OUT8_Mp9@2677_g N_VDD_Mp9@2677_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2676 N_OUT9_Mp9@2676_d N_OUT8_Mp9@2676_g N_VDD_Mp9@2676_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2675 N_OUT9_Mn9@2675_d N_OUT8_Mn9@2675_g N_VSS_Mn9@2675_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2674 N_OUT9_Mn9@2674_d N_OUT8_Mn9@2674_g N_VSS_Mn9@2674_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2675 N_OUT9_Mp9@2675_d N_OUT8_Mp9@2675_g N_VDD_Mp9@2675_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2674 N_OUT9_Mp9@2674_d N_OUT8_Mp9@2674_g N_VDD_Mp9@2674_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2673 N_OUT9_Mn9@2673_d N_OUT8_Mn9@2673_g N_VSS_Mn9@2673_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2672 N_OUT9_Mn9@2672_d N_OUT8_Mn9@2672_g N_VSS_Mn9@2672_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2673 N_OUT9_Mp9@2673_d N_OUT8_Mp9@2673_g N_VDD_Mp9@2673_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2672 N_OUT9_Mp9@2672_d N_OUT8_Mp9@2672_g N_VDD_Mp9@2672_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2671 N_OUT9_Mn9@2671_d N_OUT8_Mn9@2671_g N_VSS_Mn9@2671_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2670 N_OUT9_Mn9@2670_d N_OUT8_Mn9@2670_g N_VSS_Mn9@2670_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2671 N_OUT9_Mp9@2671_d N_OUT8_Mp9@2671_g N_VDD_Mp9@2671_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2670 N_OUT9_Mp9@2670_d N_OUT8_Mp9@2670_g N_VDD_Mp9@2670_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2669 N_OUT9_Mn9@2669_d N_OUT8_Mn9@2669_g N_VSS_Mn9@2669_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2668 N_OUT9_Mn9@2668_d N_OUT8_Mn9@2668_g N_VSS_Mn9@2668_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2669 N_OUT9_Mp9@2669_d N_OUT8_Mp9@2669_g N_VDD_Mp9@2669_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2668 N_OUT9_Mp9@2668_d N_OUT8_Mp9@2668_g N_VDD_Mp9@2668_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2667 N_OUT9_Mn9@2667_d N_OUT8_Mn9@2667_g N_VSS_Mn9@2667_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2666 N_OUT9_Mn9@2666_d N_OUT8_Mn9@2666_g N_VSS_Mn9@2666_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2667 N_OUT9_Mp9@2667_d N_OUT8_Mp9@2667_g N_VDD_Mp9@2667_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2666 N_OUT9_Mp9@2666_d N_OUT8_Mp9@2666_g N_VDD_Mp9@2666_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2665 N_OUT9_Mn9@2665_d N_OUT8_Mn9@2665_g N_VSS_Mn9@2665_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2664 N_OUT9_Mn9@2664_d N_OUT8_Mn9@2664_g N_VSS_Mn9@2664_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2665 N_OUT9_Mp9@2665_d N_OUT8_Mp9@2665_g N_VDD_Mp9@2665_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2664 N_OUT9_Mp9@2664_d N_OUT8_Mp9@2664_g N_VDD_Mp9@2664_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2663 N_OUT9_Mn9@2663_d N_OUT8_Mn9@2663_g N_VSS_Mn9@2663_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2662 N_OUT9_Mn9@2662_d N_OUT8_Mn9@2662_g N_VSS_Mn9@2662_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2663 N_OUT9_Mp9@2663_d N_OUT8_Mp9@2663_g N_VDD_Mp9@2663_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2662 N_OUT9_Mp9@2662_d N_OUT8_Mp9@2662_g N_VDD_Mp9@2662_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2661 N_OUT9_Mn9@2661_d N_OUT8_Mn9@2661_g N_VSS_Mn9@2661_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2660 N_OUT9_Mn9@2660_d N_OUT8_Mn9@2660_g N_VSS_Mn9@2660_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2661 N_OUT9_Mp9@2661_d N_OUT8_Mp9@2661_g N_VDD_Mp9@2661_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2660 N_OUT9_Mp9@2660_d N_OUT8_Mp9@2660_g N_VDD_Mp9@2660_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2659 N_OUT9_Mn9@2659_d N_OUT8_Mn9@2659_g N_VSS_Mn9@2659_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2658 N_OUT9_Mn9@2658_d N_OUT8_Mn9@2658_g N_VSS_Mn9@2658_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2659 N_OUT9_Mp9@2659_d N_OUT8_Mp9@2659_g N_VDD_Mp9@2659_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2658 N_OUT9_Mp9@2658_d N_OUT8_Mp9@2658_g N_VDD_Mp9@2658_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2657 N_OUT9_Mn9@2657_d N_OUT8_Mn9@2657_g N_VSS_Mn9@2657_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2656 N_OUT9_Mn9@2656_d N_OUT8_Mn9@2656_g N_VSS_Mn9@2656_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2657 N_OUT9_Mp9@2657_d N_OUT8_Mp9@2657_g N_VDD_Mp9@2657_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2656 N_OUT9_Mp9@2656_d N_OUT8_Mp9@2656_g N_VDD_Mp9@2656_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2655 N_OUT9_Mn9@2655_d N_OUT8_Mn9@2655_g N_VSS_Mn9@2655_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2654 N_OUT9_Mn9@2654_d N_OUT8_Mn9@2654_g N_VSS_Mn9@2654_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2655 N_OUT9_Mp9@2655_d N_OUT8_Mp9@2655_g N_VDD_Mp9@2655_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2654 N_OUT9_Mp9@2654_d N_OUT8_Mp9@2654_g N_VDD_Mp9@2654_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2653 N_OUT9_Mn9@2653_d N_OUT8_Mn9@2653_g N_VSS_Mn9@2653_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2652 N_OUT9_Mn9@2652_d N_OUT8_Mn9@2652_g N_VSS_Mn9@2652_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2653 N_OUT9_Mp9@2653_d N_OUT8_Mp9@2653_g N_VDD_Mp9@2653_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2652 N_OUT9_Mp9@2652_d N_OUT8_Mp9@2652_g N_VDD_Mp9@2652_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2651 N_OUT9_Mn9@2651_d N_OUT8_Mn9@2651_g N_VSS_Mn9@2651_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2650 N_OUT9_Mn9@2650_d N_OUT8_Mn9@2650_g N_VSS_Mn9@2650_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2651 N_OUT9_Mp9@2651_d N_OUT8_Mp9@2651_g N_VDD_Mp9@2651_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2650 N_OUT9_Mp9@2650_d N_OUT8_Mp9@2650_g N_VDD_Mp9@2650_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2649 N_OUT9_Mn9@2649_d N_OUT8_Mn9@2649_g N_VSS_Mn9@2649_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2648 N_OUT9_Mn9@2648_d N_OUT8_Mn9@2648_g N_VSS_Mn9@2648_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2649 N_OUT9_Mp9@2649_d N_OUT8_Mp9@2649_g N_VDD_Mp9@2649_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2648 N_OUT9_Mp9@2648_d N_OUT8_Mp9@2648_g N_VDD_Mp9@2648_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2647 N_OUT9_Mn9@2647_d N_OUT8_Mn9@2647_g N_VSS_Mn9@2647_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2646 N_OUT9_Mn9@2646_d N_OUT8_Mn9@2646_g N_VSS_Mn9@2646_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2647 N_OUT9_Mp9@2647_d N_OUT8_Mp9@2647_g N_VDD_Mp9@2647_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2646 N_OUT9_Mp9@2646_d N_OUT8_Mp9@2646_g N_VDD_Mp9@2646_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2645 N_OUT9_Mn9@2645_d N_OUT8_Mn9@2645_g N_VSS_Mn9@2645_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2644 N_OUT9_Mn9@2644_d N_OUT8_Mn9@2644_g N_VSS_Mn9@2644_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2645 N_OUT9_Mp9@2645_d N_OUT8_Mp9@2645_g N_VDD_Mp9@2645_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2644 N_OUT9_Mp9@2644_d N_OUT8_Mp9@2644_g N_VDD_Mp9@2644_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2643 N_OUT9_Mn9@2643_d N_OUT8_Mn9@2643_g N_VSS_Mn9@2643_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2642 N_OUT9_Mn9@2642_d N_OUT8_Mn9@2642_g N_VSS_Mn9@2642_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2643 N_OUT9_Mp9@2643_d N_OUT8_Mp9@2643_g N_VDD_Mp9@2643_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2642 N_OUT9_Mp9@2642_d N_OUT8_Mp9@2642_g N_VDD_Mp9@2642_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2641 N_OUT9_Mn9@2641_d N_OUT8_Mn9@2641_g N_VSS_Mn9@2641_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2640 N_OUT9_Mn9@2640_d N_OUT8_Mn9@2640_g N_VSS_Mn9@2640_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2641 N_OUT9_Mp9@2641_d N_OUT8_Mp9@2641_g N_VDD_Mp9@2641_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2640 N_OUT9_Mp9@2640_d N_OUT8_Mp9@2640_g N_VDD_Mp9@2640_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2639 N_OUT9_Mn9@2639_d N_OUT8_Mn9@2639_g N_VSS_Mn9@2639_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2638 N_OUT9_Mn9@2638_d N_OUT8_Mn9@2638_g N_VSS_Mn9@2638_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2639 N_OUT9_Mp9@2639_d N_OUT8_Mp9@2639_g N_VDD_Mp9@2639_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2638 N_OUT9_Mp9@2638_d N_OUT8_Mp9@2638_g N_VDD_Mp9@2638_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2637 N_OUT9_Mn9@2637_d N_OUT8_Mn9@2637_g N_VSS_Mn9@2637_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2636 N_OUT9_Mn9@2636_d N_OUT8_Mn9@2636_g N_VSS_Mn9@2636_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2637 N_OUT9_Mp9@2637_d N_OUT8_Mp9@2637_g N_VDD_Mp9@2637_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2636 N_OUT9_Mp9@2636_d N_OUT8_Mp9@2636_g N_VDD_Mp9@2636_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2635 N_OUT9_Mn9@2635_d N_OUT8_Mn9@2635_g N_VSS_Mn9@2635_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2634 N_OUT9_Mn9@2634_d N_OUT8_Mn9@2634_g N_VSS_Mn9@2634_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2635 N_OUT9_Mp9@2635_d N_OUT8_Mp9@2635_g N_VDD_Mp9@2635_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2634 N_OUT9_Mp9@2634_d N_OUT8_Mp9@2634_g N_VDD_Mp9@2634_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2633 N_OUT9_Mn9@2633_d N_OUT8_Mn9@2633_g N_VSS_Mn9@2633_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2632 N_OUT9_Mn9@2632_d N_OUT8_Mn9@2632_g N_VSS_Mn9@2632_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2633 N_OUT9_Mp9@2633_d N_OUT8_Mp9@2633_g N_VDD_Mp9@2633_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2632 N_OUT9_Mp9@2632_d N_OUT8_Mp9@2632_g N_VDD_Mp9@2632_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2631 N_OUT9_Mn9@2631_d N_OUT8_Mn9@2631_g N_VSS_Mn9@2631_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2630 N_OUT9_Mn9@2630_d N_OUT8_Mn9@2630_g N_VSS_Mn9@2630_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2631 N_OUT9_Mp9@2631_d N_OUT8_Mp9@2631_g N_VDD_Mp9@2631_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2630 N_OUT9_Mp9@2630_d N_OUT8_Mp9@2630_g N_VDD_Mp9@2630_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2629 N_OUT9_Mn9@2629_d N_OUT8_Mn9@2629_g N_VSS_Mn9@2629_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2628 N_OUT9_Mn9@2628_d N_OUT8_Mn9@2628_g N_VSS_Mn9@2628_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2629 N_OUT9_Mp9@2629_d N_OUT8_Mp9@2629_g N_VDD_Mp9@2629_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2628 N_OUT9_Mp9@2628_d N_OUT8_Mp9@2628_g N_VDD_Mp9@2628_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2627 N_OUT9_Mn9@2627_d N_OUT8_Mn9@2627_g N_VSS_Mn9@2627_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2626 N_OUT9_Mn9@2626_d N_OUT8_Mn9@2626_g N_VSS_Mn9@2626_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2627 N_OUT9_Mp9@2627_d N_OUT8_Mp9@2627_g N_VDD_Mp9@2627_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2626 N_OUT9_Mp9@2626_d N_OUT8_Mp9@2626_g N_VDD_Mp9@2626_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2625 N_OUT9_Mn9@2625_d N_OUT8_Mn9@2625_g N_VSS_Mn9@2625_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2624 N_OUT9_Mn9@2624_d N_OUT8_Mn9@2624_g N_VSS_Mn9@2624_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2625 N_OUT9_Mp9@2625_d N_OUT8_Mp9@2625_g N_VDD_Mp9@2625_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2624 N_OUT9_Mp9@2624_d N_OUT8_Mp9@2624_g N_VDD_Mp9@2624_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2623 N_OUT9_Mn9@2623_d N_OUT8_Mn9@2623_g N_VSS_Mn9@2623_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2622 N_OUT9_Mn9@2622_d N_OUT8_Mn9@2622_g N_VSS_Mn9@2622_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2623 N_OUT9_Mp9@2623_d N_OUT8_Mp9@2623_g N_VDD_Mp9@2623_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2622 N_OUT9_Mp9@2622_d N_OUT8_Mp9@2622_g N_VDD_Mp9@2622_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2621 N_OUT9_Mn9@2621_d N_OUT8_Mn9@2621_g N_VSS_Mn9@2621_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2620 N_OUT9_Mn9@2620_d N_OUT8_Mn9@2620_g N_VSS_Mn9@2620_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2621 N_OUT9_Mp9@2621_d N_OUT8_Mp9@2621_g N_VDD_Mp9@2621_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2620 N_OUT9_Mp9@2620_d N_OUT8_Mp9@2620_g N_VDD_Mp9@2620_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2619 N_OUT9_Mn9@2619_d N_OUT8_Mn9@2619_g N_VSS_Mn9@2619_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2618 N_OUT9_Mn9@2618_d N_OUT8_Mn9@2618_g N_VSS_Mn9@2618_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2619 N_OUT9_Mp9@2619_d N_OUT8_Mp9@2619_g N_VDD_Mp9@2619_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2618 N_OUT9_Mp9@2618_d N_OUT8_Mp9@2618_g N_VDD_Mp9@2618_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2617 N_OUT9_Mn9@2617_d N_OUT8_Mn9@2617_g N_VSS_Mn9@2617_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2616 N_OUT9_Mn9@2616_d N_OUT8_Mn9@2616_g N_VSS_Mn9@2616_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2617 N_OUT9_Mp9@2617_d N_OUT8_Mp9@2617_g N_VDD_Mp9@2617_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2616 N_OUT9_Mp9@2616_d N_OUT8_Mp9@2616_g N_VDD_Mp9@2616_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2615 N_OUT9_Mn9@2615_d N_OUT8_Mn9@2615_g N_VSS_Mn9@2615_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2614 N_OUT9_Mn9@2614_d N_OUT8_Mn9@2614_g N_VSS_Mn9@2614_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2615 N_OUT9_Mp9@2615_d N_OUT8_Mp9@2615_g N_VDD_Mp9@2615_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2614 N_OUT9_Mp9@2614_d N_OUT8_Mp9@2614_g N_VDD_Mp9@2614_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2613 N_OUT9_Mn9@2613_d N_OUT8_Mn9@2613_g N_VSS_Mn9@2613_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2612 N_OUT9_Mn9@2612_d N_OUT8_Mn9@2612_g N_VSS_Mn9@2612_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2613 N_OUT9_Mp9@2613_d N_OUT8_Mp9@2613_g N_VDD_Mp9@2613_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2612 N_OUT9_Mp9@2612_d N_OUT8_Mp9@2612_g N_VDD_Mp9@2612_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2611 N_OUT9_Mn9@2611_d N_OUT8_Mn9@2611_g N_VSS_Mn9@2611_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2610 N_OUT9_Mn9@2610_d N_OUT8_Mn9@2610_g N_VSS_Mn9@2610_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2611 N_OUT9_Mp9@2611_d N_OUT8_Mp9@2611_g N_VDD_Mp9@2611_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2610 N_OUT9_Mp9@2610_d N_OUT8_Mp9@2610_g N_VDD_Mp9@2610_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2609 N_OUT9_Mn9@2609_d N_OUT8_Mn9@2609_g N_VSS_Mn9@2609_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2608 N_OUT9_Mn9@2608_d N_OUT8_Mn9@2608_g N_VSS_Mn9@2608_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2609 N_OUT9_Mp9@2609_d N_OUT8_Mp9@2609_g N_VDD_Mp9@2609_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2608 N_OUT9_Mp9@2608_d N_OUT8_Mp9@2608_g N_VDD_Mp9@2608_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2607 N_OUT9_Mn9@2607_d N_OUT8_Mn9@2607_g N_VSS_Mn9@2607_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2606 N_OUT9_Mn9@2606_d N_OUT8_Mn9@2606_g N_VSS_Mn9@2606_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2607 N_OUT9_Mp9@2607_d N_OUT8_Mp9@2607_g N_VDD_Mp9@2607_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2606 N_OUT9_Mp9@2606_d N_OUT8_Mp9@2606_g N_VDD_Mp9@2606_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2605 N_OUT9_Mn9@2605_d N_OUT8_Mn9@2605_g N_VSS_Mn9@2605_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2604 N_OUT9_Mn9@2604_d N_OUT8_Mn9@2604_g N_VSS_Mn9@2604_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2605 N_OUT9_Mp9@2605_d N_OUT8_Mp9@2605_g N_VDD_Mp9@2605_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2604 N_OUT9_Mp9@2604_d N_OUT8_Mp9@2604_g N_VDD_Mp9@2604_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2603 N_OUT9_Mn9@2603_d N_OUT8_Mn9@2603_g N_VSS_Mn9@2603_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2602 N_OUT9_Mn9@2602_d N_OUT8_Mn9@2602_g N_VSS_Mn9@2602_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2603 N_OUT9_Mp9@2603_d N_OUT8_Mp9@2603_g N_VDD_Mp9@2603_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2602 N_OUT9_Mp9@2602_d N_OUT8_Mp9@2602_g N_VDD_Mp9@2602_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2601 N_OUT9_Mn9@2601_d N_OUT8_Mn9@2601_g N_VSS_Mn9@2601_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2600 N_OUT9_Mn9@2600_d N_OUT8_Mn9@2600_g N_VSS_Mn9@2600_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2601 N_OUT9_Mp9@2601_d N_OUT8_Mp9@2601_g N_VDD_Mp9@2601_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2600 N_OUT9_Mp9@2600_d N_OUT8_Mp9@2600_g N_VDD_Mp9@2600_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2599 N_OUT9_Mn9@2599_d N_OUT8_Mn9@2599_g N_VSS_Mn9@2599_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2598 N_OUT9_Mn9@2598_d N_OUT8_Mn9@2598_g N_VSS_Mn9@2598_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2599 N_OUT9_Mp9@2599_d N_OUT8_Mp9@2599_g N_VDD_Mp9@2599_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2598 N_OUT9_Mp9@2598_d N_OUT8_Mp9@2598_g N_VDD_Mp9@2598_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2597 N_OUT9_Mn9@2597_d N_OUT8_Mn9@2597_g N_VSS_Mn9@2597_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2596 N_OUT9_Mn9@2596_d N_OUT8_Mn9@2596_g N_VSS_Mn9@2596_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2597 N_OUT9_Mp9@2597_d N_OUT8_Mp9@2597_g N_VDD_Mp9@2597_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2596 N_OUT9_Mp9@2596_d N_OUT8_Mp9@2596_g N_VDD_Mp9@2596_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2595 N_OUT9_Mn9@2595_d N_OUT8_Mn9@2595_g N_VSS_Mn9@2595_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2594 N_OUT9_Mn9@2594_d N_OUT8_Mn9@2594_g N_VSS_Mn9@2594_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2595 N_OUT9_Mp9@2595_d N_OUT8_Mp9@2595_g N_VDD_Mp9@2595_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2594 N_OUT9_Mp9@2594_d N_OUT8_Mp9@2594_g N_VDD_Mp9@2594_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2593 N_OUT9_Mn9@2593_d N_OUT8_Mn9@2593_g N_VSS_Mn9@2593_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2592 N_OUT9_Mn9@2592_d N_OUT8_Mn9@2592_g N_VSS_Mn9@2592_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2593 N_OUT9_Mp9@2593_d N_OUT8_Mp9@2593_g N_VDD_Mp9@2593_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2592 N_OUT9_Mp9@2592_d N_OUT8_Mp9@2592_g N_VDD_Mp9@2592_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2591 N_OUT9_Mn9@2591_d N_OUT8_Mn9@2591_g N_VSS_Mn9@2591_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2590 N_OUT9_Mn9@2590_d N_OUT8_Mn9@2590_g N_VSS_Mn9@2590_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2591 N_OUT9_Mp9@2591_d N_OUT8_Mp9@2591_g N_VDD_Mp9@2591_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2590 N_OUT9_Mp9@2590_d N_OUT8_Mp9@2590_g N_VDD_Mp9@2590_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2589 N_OUT9_Mn9@2589_d N_OUT8_Mn9@2589_g N_VSS_Mn9@2589_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2588 N_OUT9_Mn9@2588_d N_OUT8_Mn9@2588_g N_VSS_Mn9@2588_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2589 N_OUT9_Mp9@2589_d N_OUT8_Mp9@2589_g N_VDD_Mp9@2589_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2588 N_OUT9_Mp9@2588_d N_OUT8_Mp9@2588_g N_VDD_Mp9@2588_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2587 N_OUT9_Mn9@2587_d N_OUT8_Mn9@2587_g N_VSS_Mn9@2587_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2586 N_OUT9_Mn9@2586_d N_OUT8_Mn9@2586_g N_VSS_Mn9@2586_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2587 N_OUT9_Mp9@2587_d N_OUT8_Mp9@2587_g N_VDD_Mp9@2587_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2586 N_OUT9_Mp9@2586_d N_OUT8_Mp9@2586_g N_VDD_Mp9@2586_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2585 N_OUT9_Mn9@2585_d N_OUT8_Mn9@2585_g N_VSS_Mn9@2585_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2584 N_OUT9_Mn9@2584_d N_OUT8_Mn9@2584_g N_VSS_Mn9@2584_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2585 N_OUT9_Mp9@2585_d N_OUT8_Mp9@2585_g N_VDD_Mp9@2585_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2584 N_OUT9_Mp9@2584_d N_OUT8_Mp9@2584_g N_VDD_Mp9@2584_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2583 N_OUT9_Mn9@2583_d N_OUT8_Mn9@2583_g N_VSS_Mn9@2583_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2582 N_OUT9_Mn9@2582_d N_OUT8_Mn9@2582_g N_VSS_Mn9@2582_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2583 N_OUT9_Mp9@2583_d N_OUT8_Mp9@2583_g N_VDD_Mp9@2583_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2582 N_OUT9_Mp9@2582_d N_OUT8_Mp9@2582_g N_VDD_Mp9@2582_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2581 N_OUT9_Mn9@2581_d N_OUT8_Mn9@2581_g N_VSS_Mn9@2581_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2580 N_OUT9_Mn9@2580_d N_OUT8_Mn9@2580_g N_VSS_Mn9@2580_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2581 N_OUT9_Mp9@2581_d N_OUT8_Mp9@2581_g N_VDD_Mp9@2581_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2580 N_OUT9_Mp9@2580_d N_OUT8_Mp9@2580_g N_VDD_Mp9@2580_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2579 N_OUT9_Mn9@2579_d N_OUT8_Mn9@2579_g N_VSS_Mn9@2579_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2578 N_OUT9_Mn9@2578_d N_OUT8_Mn9@2578_g N_VSS_Mn9@2578_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2579 N_OUT9_Mp9@2579_d N_OUT8_Mp9@2579_g N_VDD_Mp9@2579_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2578 N_OUT9_Mp9@2578_d N_OUT8_Mp9@2578_g N_VDD_Mp9@2578_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2577 N_OUT9_Mn9@2577_d N_OUT8_Mn9@2577_g N_VSS_Mn9@2577_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2576 N_OUT9_Mn9@2576_d N_OUT8_Mn9@2576_g N_VSS_Mn9@2576_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2577 N_OUT9_Mp9@2577_d N_OUT8_Mp9@2577_g N_VDD_Mp9@2577_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2576 N_OUT9_Mp9@2576_d N_OUT8_Mp9@2576_g N_VDD_Mp9@2576_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2575 N_OUT9_Mn9@2575_d N_OUT8_Mn9@2575_g N_VSS_Mn9@2575_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2574 N_OUT9_Mn9@2574_d N_OUT8_Mn9@2574_g N_VSS_Mn9@2574_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2575 N_OUT9_Mp9@2575_d N_OUT8_Mp9@2575_g N_VDD_Mp9@2575_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2574 N_OUT9_Mp9@2574_d N_OUT8_Mp9@2574_g N_VDD_Mp9@2574_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2573 N_OUT9_Mn9@2573_d N_OUT8_Mn9@2573_g N_VSS_Mn9@2573_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2572 N_OUT9_Mn9@2572_d N_OUT8_Mn9@2572_g N_VSS_Mn9@2572_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2573 N_OUT9_Mp9@2573_d N_OUT8_Mp9@2573_g N_VDD_Mp9@2573_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2572 N_OUT9_Mp9@2572_d N_OUT8_Mp9@2572_g N_VDD_Mp9@2572_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2571 N_OUT9_Mn9@2571_d N_OUT8_Mn9@2571_g N_VSS_Mn9@2571_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2570 N_OUT9_Mn9@2570_d N_OUT8_Mn9@2570_g N_VSS_Mn9@2570_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2571 N_OUT9_Mp9@2571_d N_OUT8_Mp9@2571_g N_VDD_Mp9@2571_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2570 N_OUT9_Mp9@2570_d N_OUT8_Mp9@2570_g N_VDD_Mp9@2570_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2569 N_OUT9_Mn9@2569_d N_OUT8_Mn9@2569_g N_VSS_Mn9@2569_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2568 N_OUT9_Mn9@2568_d N_OUT8_Mn9@2568_g N_VSS_Mn9@2568_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2569 N_OUT9_Mp9@2569_d N_OUT8_Mp9@2569_g N_VDD_Mp9@2569_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2568 N_OUT9_Mp9@2568_d N_OUT8_Mp9@2568_g N_VDD_Mp9@2568_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2567 N_OUT9_Mn9@2567_d N_OUT8_Mn9@2567_g N_VSS_Mn9@2567_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2566 N_OUT9_Mn9@2566_d N_OUT8_Mn9@2566_g N_VSS_Mn9@2566_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2567 N_OUT9_Mp9@2567_d N_OUT8_Mp9@2567_g N_VDD_Mp9@2567_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2566 N_OUT9_Mp9@2566_d N_OUT8_Mp9@2566_g N_VDD_Mp9@2566_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2565 N_OUT9_Mn9@2565_d N_OUT8_Mn9@2565_g N_VSS_Mn9@2565_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2564 N_OUT9_Mn9@2564_d N_OUT8_Mn9@2564_g N_VSS_Mn9@2564_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2565 N_OUT9_Mp9@2565_d N_OUT8_Mp9@2565_g N_VDD_Mp9@2565_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2564 N_OUT9_Mp9@2564_d N_OUT8_Mp9@2564_g N_VDD_Mp9@2564_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2563 N_OUT9_Mn9@2563_d N_OUT8_Mn9@2563_g N_VSS_Mn9@2563_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2562 N_OUT9_Mn9@2562_d N_OUT8_Mn9@2562_g N_VSS_Mn9@2562_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2563 N_OUT9_Mp9@2563_d N_OUT8_Mp9@2563_g N_VDD_Mp9@2563_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2562 N_OUT9_Mp9@2562_d N_OUT8_Mp9@2562_g N_VDD_Mp9@2562_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2561 N_OUT9_Mn9@2561_d N_OUT8_Mn9@2561_g N_VSS_Mn9@2561_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2560 N_OUT9_Mn9@2560_d N_OUT8_Mn9@2560_g N_VSS_Mn9@2560_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2561 N_OUT9_Mp9@2561_d N_OUT8_Mp9@2561_g N_VDD_Mp9@2561_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2560 N_OUT9_Mp9@2560_d N_OUT8_Mp9@2560_g N_VDD_Mp9@2560_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2559 N_OUT9_Mn9@2559_d N_OUT8_Mn9@2559_g N_VSS_Mn9@2559_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2558 N_OUT9_Mn9@2558_d N_OUT8_Mn9@2558_g N_VSS_Mn9@2558_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2559 N_OUT9_Mp9@2559_d N_OUT8_Mp9@2559_g N_VDD_Mp9@2559_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2558 N_OUT9_Mp9@2558_d N_OUT8_Mp9@2558_g N_VDD_Mp9@2558_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2557 N_OUT9_Mn9@2557_d N_OUT8_Mn9@2557_g N_VSS_Mn9@2557_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2556 N_OUT9_Mn9@2556_d N_OUT8_Mn9@2556_g N_VSS_Mn9@2556_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2557 N_OUT9_Mp9@2557_d N_OUT8_Mp9@2557_g N_VDD_Mp9@2557_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2556 N_OUT9_Mp9@2556_d N_OUT8_Mp9@2556_g N_VDD_Mp9@2556_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2555 N_OUT9_Mn9@2555_d N_OUT8_Mn9@2555_g N_VSS_Mn9@2555_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2554 N_OUT9_Mn9@2554_d N_OUT8_Mn9@2554_g N_VSS_Mn9@2554_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2555 N_OUT9_Mp9@2555_d N_OUT8_Mp9@2555_g N_VDD_Mp9@2555_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2554 N_OUT9_Mp9@2554_d N_OUT8_Mp9@2554_g N_VDD_Mp9@2554_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2553 N_OUT9_Mn9@2553_d N_OUT8_Mn9@2553_g N_VSS_Mn9@2553_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2552 N_OUT9_Mn9@2552_d N_OUT8_Mn9@2552_g N_VSS_Mn9@2552_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2553 N_OUT9_Mp9@2553_d N_OUT8_Mp9@2553_g N_VDD_Mp9@2553_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2552 N_OUT9_Mp9@2552_d N_OUT8_Mp9@2552_g N_VDD_Mp9@2552_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2551 N_OUT9_Mn9@2551_d N_OUT8_Mn9@2551_g N_VSS_Mn9@2551_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2550 N_OUT9_Mn9@2550_d N_OUT8_Mn9@2550_g N_VSS_Mn9@2550_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2551 N_OUT9_Mp9@2551_d N_OUT8_Mp9@2551_g N_VDD_Mp9@2551_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2550 N_OUT9_Mp9@2550_d N_OUT8_Mp9@2550_g N_VDD_Mp9@2550_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2549 N_OUT9_Mn9@2549_d N_OUT8_Mn9@2549_g N_VSS_Mn9@2549_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2548 N_OUT9_Mn9@2548_d N_OUT8_Mn9@2548_g N_VSS_Mn9@2548_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2549 N_OUT9_Mp9@2549_d N_OUT8_Mp9@2549_g N_VDD_Mp9@2549_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2548 N_OUT9_Mp9@2548_d N_OUT8_Mp9@2548_g N_VDD_Mp9@2548_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2547 N_OUT9_Mn9@2547_d N_OUT8_Mn9@2547_g N_VSS_Mn9@2547_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2546 N_OUT9_Mn9@2546_d N_OUT8_Mn9@2546_g N_VSS_Mn9@2546_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2547 N_OUT9_Mp9@2547_d N_OUT8_Mp9@2547_g N_VDD_Mp9@2547_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2546 N_OUT9_Mp9@2546_d N_OUT8_Mp9@2546_g N_VDD_Mp9@2546_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2545 N_OUT9_Mn9@2545_d N_OUT8_Mn9@2545_g N_VSS_Mn9@2545_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2544 N_OUT9_Mn9@2544_d N_OUT8_Mn9@2544_g N_VSS_Mn9@2544_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2545 N_OUT9_Mp9@2545_d N_OUT8_Mp9@2545_g N_VDD_Mp9@2545_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2544 N_OUT9_Mp9@2544_d N_OUT8_Mp9@2544_g N_VDD_Mp9@2544_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2543 N_OUT9_Mn9@2543_d N_OUT8_Mn9@2543_g N_VSS_Mn9@2543_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2542 N_OUT9_Mn9@2542_d N_OUT8_Mn9@2542_g N_VSS_Mn9@2542_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2543 N_OUT9_Mp9@2543_d N_OUT8_Mp9@2543_g N_VDD_Mp9@2543_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2542 N_OUT9_Mp9@2542_d N_OUT8_Mp9@2542_g N_VDD_Mp9@2542_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2541 N_OUT9_Mn9@2541_d N_OUT8_Mn9@2541_g N_VSS_Mn9@2541_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2540 N_OUT9_Mn9@2540_d N_OUT8_Mn9@2540_g N_VSS_Mn9@2540_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2541 N_OUT9_Mp9@2541_d N_OUT8_Mp9@2541_g N_VDD_Mp9@2541_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2540 N_OUT9_Mp9@2540_d N_OUT8_Mp9@2540_g N_VDD_Mp9@2540_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2539 N_OUT9_Mn9@2539_d N_OUT8_Mn9@2539_g N_VSS_Mn9@2539_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2538 N_OUT9_Mn9@2538_d N_OUT8_Mn9@2538_g N_VSS_Mn9@2538_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2539 N_OUT9_Mp9@2539_d N_OUT8_Mp9@2539_g N_VDD_Mp9@2539_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2538 N_OUT9_Mp9@2538_d N_OUT8_Mp9@2538_g N_VDD_Mp9@2538_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2537 N_OUT9_Mn9@2537_d N_OUT8_Mn9@2537_g N_VSS_Mn9@2537_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2536 N_OUT9_Mn9@2536_d N_OUT8_Mn9@2536_g N_VSS_Mn9@2536_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2537 N_OUT9_Mp9@2537_d N_OUT8_Mp9@2537_g N_VDD_Mp9@2537_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2536 N_OUT9_Mp9@2536_d N_OUT8_Mp9@2536_g N_VDD_Mp9@2536_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2535 N_OUT9_Mn9@2535_d N_OUT8_Mn9@2535_g N_VSS_Mn9@2535_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2534 N_OUT9_Mn9@2534_d N_OUT8_Mn9@2534_g N_VSS_Mn9@2534_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2535 N_OUT9_Mp9@2535_d N_OUT8_Mp9@2535_g N_VDD_Mp9@2535_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2534 N_OUT9_Mp9@2534_d N_OUT8_Mp9@2534_g N_VDD_Mp9@2534_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2533 N_OUT9_Mn9@2533_d N_OUT8_Mn9@2533_g N_VSS_Mn9@2533_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2532 N_OUT9_Mn9@2532_d N_OUT8_Mn9@2532_g N_VSS_Mn9@2532_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2533 N_OUT9_Mp9@2533_d N_OUT8_Mp9@2533_g N_VDD_Mp9@2533_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2532 N_OUT9_Mp9@2532_d N_OUT8_Mp9@2532_g N_VDD_Mp9@2532_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2531 N_OUT9_Mn9@2531_d N_OUT8_Mn9@2531_g N_VSS_Mn9@2531_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2530 N_OUT9_Mn9@2530_d N_OUT8_Mn9@2530_g N_VSS_Mn9@2530_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2531 N_OUT9_Mp9@2531_d N_OUT8_Mp9@2531_g N_VDD_Mp9@2531_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2530 N_OUT9_Mp9@2530_d N_OUT8_Mp9@2530_g N_VDD_Mp9@2530_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2529 N_OUT9_Mn9@2529_d N_OUT8_Mn9@2529_g N_VSS_Mn9@2529_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2528 N_OUT9_Mn9@2528_d N_OUT8_Mn9@2528_g N_VSS_Mn9@2528_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2529 N_OUT9_Mp9@2529_d N_OUT8_Mp9@2529_g N_VDD_Mp9@2529_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2528 N_OUT9_Mp9@2528_d N_OUT8_Mp9@2528_g N_VDD_Mp9@2528_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2527 N_OUT9_Mn9@2527_d N_OUT8_Mn9@2527_g N_VSS_Mn9@2527_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2526 N_OUT9_Mn9@2526_d N_OUT8_Mn9@2526_g N_VSS_Mn9@2526_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2527 N_OUT9_Mp9@2527_d N_OUT8_Mp9@2527_g N_VDD_Mp9@2527_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2526 N_OUT9_Mp9@2526_d N_OUT8_Mp9@2526_g N_VDD_Mp9@2526_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2525 N_OUT9_Mn9@2525_d N_OUT8_Mn9@2525_g N_VSS_Mn9@2525_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2524 N_OUT9_Mn9@2524_d N_OUT8_Mn9@2524_g N_VSS_Mn9@2524_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2525 N_OUT9_Mp9@2525_d N_OUT8_Mp9@2525_g N_VDD_Mp9@2525_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2524 N_OUT9_Mp9@2524_d N_OUT8_Mp9@2524_g N_VDD_Mp9@2524_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2523 N_OUT9_Mn9@2523_d N_OUT8_Mn9@2523_g N_VSS_Mn9@2523_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2522 N_OUT9_Mn9@2522_d N_OUT8_Mn9@2522_g N_VSS_Mn9@2522_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2523 N_OUT9_Mp9@2523_d N_OUT8_Mp9@2523_g N_VDD_Mp9@2523_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2522 N_OUT9_Mp9@2522_d N_OUT8_Mp9@2522_g N_VDD_Mp9@2522_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2521 N_OUT9_Mn9@2521_d N_OUT8_Mn9@2521_g N_VSS_Mn9@2521_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2520 N_OUT9_Mn9@2520_d N_OUT8_Mn9@2520_g N_VSS_Mn9@2520_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2521 N_OUT9_Mp9@2521_d N_OUT8_Mp9@2521_g N_VDD_Mp9@2521_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2520 N_OUT9_Mp9@2520_d N_OUT8_Mp9@2520_g N_VDD_Mp9@2520_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2519 N_OUT9_Mn9@2519_d N_OUT8_Mn9@2519_g N_VSS_Mn9@2519_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2518 N_OUT9_Mn9@2518_d N_OUT8_Mn9@2518_g N_VSS_Mn9@2518_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2519 N_OUT9_Mp9@2519_d N_OUT8_Mp9@2519_g N_VDD_Mp9@2519_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2518 N_OUT9_Mp9@2518_d N_OUT8_Mp9@2518_g N_VDD_Mp9@2518_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2517 N_OUT9_Mn9@2517_d N_OUT8_Mn9@2517_g N_VSS_Mn9@2517_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2516 N_OUT9_Mn9@2516_d N_OUT8_Mn9@2516_g N_VSS_Mn9@2516_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2517 N_OUT9_Mp9@2517_d N_OUT8_Mp9@2517_g N_VDD_Mp9@2517_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2516 N_OUT9_Mp9@2516_d N_OUT8_Mp9@2516_g N_VDD_Mp9@2516_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2515 N_OUT9_Mn9@2515_d N_OUT8_Mn9@2515_g N_VSS_Mn9@2515_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2514 N_OUT9_Mn9@2514_d N_OUT8_Mn9@2514_g N_VSS_Mn9@2514_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2515 N_OUT9_Mp9@2515_d N_OUT8_Mp9@2515_g N_VDD_Mp9@2515_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2514 N_OUT9_Mp9@2514_d N_OUT8_Mp9@2514_g N_VDD_Mp9@2514_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2513 N_OUT9_Mn9@2513_d N_OUT8_Mn9@2513_g N_VSS_Mn9@2513_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2512 N_OUT9_Mn9@2512_d N_OUT8_Mn9@2512_g N_VSS_Mn9@2512_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2513 N_OUT9_Mp9@2513_d N_OUT8_Mp9@2513_g N_VDD_Mp9@2513_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2512 N_OUT9_Mp9@2512_d N_OUT8_Mp9@2512_g N_VDD_Mp9@2512_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2511 N_OUT9_Mn9@2511_d N_OUT8_Mn9@2511_g N_VSS_Mn9@2511_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2510 N_OUT9_Mn9@2510_d N_OUT8_Mn9@2510_g N_VSS_Mn9@2510_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2511 N_OUT9_Mp9@2511_d N_OUT8_Mp9@2511_g N_VDD_Mp9@2511_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2510 N_OUT9_Mp9@2510_d N_OUT8_Mp9@2510_g N_VDD_Mp9@2510_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2509 N_OUT9_Mn9@2509_d N_OUT8_Mn9@2509_g N_VSS_Mn9@2509_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2508 N_OUT9_Mn9@2508_d N_OUT8_Mn9@2508_g N_VSS_Mn9@2508_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2509 N_OUT9_Mp9@2509_d N_OUT8_Mp9@2509_g N_VDD_Mp9@2509_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2508 N_OUT9_Mp9@2508_d N_OUT8_Mp9@2508_g N_VDD_Mp9@2508_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2507 N_OUT9_Mn9@2507_d N_OUT8_Mn9@2507_g N_VSS_Mn9@2507_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2506 N_OUT9_Mn9@2506_d N_OUT8_Mn9@2506_g N_VSS_Mn9@2506_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2507 N_OUT9_Mp9@2507_d N_OUT8_Mp9@2507_g N_VDD_Mp9@2507_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2506 N_OUT9_Mp9@2506_d N_OUT8_Mp9@2506_g N_VDD_Mp9@2506_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2505 N_OUT9_Mn9@2505_d N_OUT8_Mn9@2505_g N_VSS_Mn9@2505_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2504 N_OUT9_Mn9@2504_d N_OUT8_Mn9@2504_g N_VSS_Mn9@2504_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2505 N_OUT9_Mp9@2505_d N_OUT8_Mp9@2505_g N_VDD_Mp9@2505_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2504 N_OUT9_Mp9@2504_d N_OUT8_Mp9@2504_g N_VDD_Mp9@2504_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2503 N_OUT9_Mn9@2503_d N_OUT8_Mn9@2503_g N_VSS_Mn9@2503_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2502 N_OUT9_Mn9@2502_d N_OUT8_Mn9@2502_g N_VSS_Mn9@2502_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2503 N_OUT9_Mp9@2503_d N_OUT8_Mp9@2503_g N_VDD_Mp9@2503_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2502 N_OUT9_Mp9@2502_d N_OUT8_Mp9@2502_g N_VDD_Mp9@2502_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2501 N_OUT9_Mn9@2501_d N_OUT8_Mn9@2501_g N_VSS_Mn9@2501_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2500 N_OUT9_Mn9@2500_d N_OUT8_Mn9@2500_g N_VSS_Mn9@2500_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2501 N_OUT9_Mp9@2501_d N_OUT8_Mp9@2501_g N_VDD_Mp9@2501_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2500 N_OUT9_Mp9@2500_d N_OUT8_Mp9@2500_g N_VDD_Mp9@2500_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2499 N_OUT9_Mn9@2499_d N_OUT8_Mn9@2499_g N_VSS_Mn9@2499_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2498 N_OUT9_Mn9@2498_d N_OUT8_Mn9@2498_g N_VSS_Mn9@2498_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2499 N_OUT9_Mp9@2499_d N_OUT8_Mp9@2499_g N_VDD_Mp9@2499_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2498 N_OUT9_Mp9@2498_d N_OUT8_Mp9@2498_g N_VDD_Mp9@2498_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2497 N_OUT9_Mn9@2497_d N_OUT8_Mn9@2497_g N_VSS_Mn9@2497_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2496 N_OUT9_Mn9@2496_d N_OUT8_Mn9@2496_g N_VSS_Mn9@2496_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2497 N_OUT9_Mp9@2497_d N_OUT8_Mp9@2497_g N_VDD_Mp9@2497_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2496 N_OUT9_Mp9@2496_d N_OUT8_Mp9@2496_g N_VDD_Mp9@2496_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2495 N_OUT9_Mn9@2495_d N_OUT8_Mn9@2495_g N_VSS_Mn9@2495_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2494 N_OUT9_Mn9@2494_d N_OUT8_Mn9@2494_g N_VSS_Mn9@2494_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2495 N_OUT9_Mp9@2495_d N_OUT8_Mp9@2495_g N_VDD_Mp9@2495_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2494 N_OUT9_Mp9@2494_d N_OUT8_Mp9@2494_g N_VDD_Mp9@2494_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2493 N_OUT9_Mn9@2493_d N_OUT8_Mn9@2493_g N_VSS_Mn9@2493_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2492 N_OUT9_Mn9@2492_d N_OUT8_Mn9@2492_g N_VSS_Mn9@2492_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2493 N_OUT9_Mp9@2493_d N_OUT8_Mp9@2493_g N_VDD_Mp9@2493_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2492 N_OUT9_Mp9@2492_d N_OUT8_Mp9@2492_g N_VDD_Mp9@2492_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2491 N_OUT9_Mn9@2491_d N_OUT8_Mn9@2491_g N_VSS_Mn9@2491_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2490 N_OUT9_Mn9@2490_d N_OUT8_Mn9@2490_g N_VSS_Mn9@2490_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2491 N_OUT9_Mp9@2491_d N_OUT8_Mp9@2491_g N_VDD_Mp9@2491_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2490 N_OUT9_Mp9@2490_d N_OUT8_Mp9@2490_g N_VDD_Mp9@2490_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2489 N_OUT9_Mn9@2489_d N_OUT8_Mn9@2489_g N_VSS_Mn9@2489_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2488 N_OUT9_Mn9@2488_d N_OUT8_Mn9@2488_g N_VSS_Mn9@2488_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2489 N_OUT9_Mp9@2489_d N_OUT8_Mp9@2489_g N_VDD_Mp9@2489_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2488 N_OUT9_Mp9@2488_d N_OUT8_Mp9@2488_g N_VDD_Mp9@2488_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2487 N_OUT9_Mn9@2487_d N_OUT8_Mn9@2487_g N_VSS_Mn9@2487_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2486 N_OUT9_Mn9@2486_d N_OUT8_Mn9@2486_g N_VSS_Mn9@2486_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2487 N_OUT9_Mp9@2487_d N_OUT8_Mp9@2487_g N_VDD_Mp9@2487_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2486 N_OUT9_Mp9@2486_d N_OUT8_Mp9@2486_g N_VDD_Mp9@2486_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2485 N_OUT9_Mn9@2485_d N_OUT8_Mn9@2485_g N_VSS_Mn9@2485_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2484 N_OUT9_Mn9@2484_d N_OUT8_Mn9@2484_g N_VSS_Mn9@2484_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2485 N_OUT9_Mp9@2485_d N_OUT8_Mp9@2485_g N_VDD_Mp9@2485_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2484 N_OUT9_Mp9@2484_d N_OUT8_Mp9@2484_g N_VDD_Mp9@2484_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2483 N_OUT9_Mn9@2483_d N_OUT8_Mn9@2483_g N_VSS_Mn9@2483_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2482 N_OUT9_Mn9@2482_d N_OUT8_Mn9@2482_g N_VSS_Mn9@2482_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2483 N_OUT9_Mp9@2483_d N_OUT8_Mp9@2483_g N_VDD_Mp9@2483_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2482 N_OUT9_Mp9@2482_d N_OUT8_Mp9@2482_g N_VDD_Mp9@2482_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2481 N_OUT9_Mn9@2481_d N_OUT8_Mn9@2481_g N_VSS_Mn9@2481_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2480 N_OUT9_Mn9@2480_d N_OUT8_Mn9@2480_g N_VSS_Mn9@2480_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2481 N_OUT9_Mp9@2481_d N_OUT8_Mp9@2481_g N_VDD_Mp9@2481_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2480 N_OUT9_Mp9@2480_d N_OUT8_Mp9@2480_g N_VDD_Mp9@2480_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2479 N_OUT9_Mn9@2479_d N_OUT8_Mn9@2479_g N_VSS_Mn9@2479_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2478 N_OUT9_Mn9@2478_d N_OUT8_Mn9@2478_g N_VSS_Mn9@2478_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2479 N_OUT9_Mp9@2479_d N_OUT8_Mp9@2479_g N_VDD_Mp9@2479_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2478 N_OUT9_Mp9@2478_d N_OUT8_Mp9@2478_g N_VDD_Mp9@2478_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2477 N_OUT9_Mn9@2477_d N_OUT8_Mn9@2477_g N_VSS_Mn9@2477_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2476 N_OUT9_Mn9@2476_d N_OUT8_Mn9@2476_g N_VSS_Mn9@2476_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2477 N_OUT9_Mp9@2477_d N_OUT8_Mp9@2477_g N_VDD_Mp9@2477_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2476 N_OUT9_Mp9@2476_d N_OUT8_Mp9@2476_g N_VDD_Mp9@2476_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2475 N_OUT9_Mn9@2475_d N_OUT8_Mn9@2475_g N_VSS_Mn9@2475_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2474 N_OUT9_Mn9@2474_d N_OUT8_Mn9@2474_g N_VSS_Mn9@2474_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2475 N_OUT9_Mp9@2475_d N_OUT8_Mp9@2475_g N_VDD_Mp9@2475_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2474 N_OUT9_Mp9@2474_d N_OUT8_Mp9@2474_g N_VDD_Mp9@2474_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2473 N_OUT9_Mn9@2473_d N_OUT8_Mn9@2473_g N_VSS_Mn9@2473_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2472 N_OUT9_Mn9@2472_d N_OUT8_Mn9@2472_g N_VSS_Mn9@2472_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2473 N_OUT9_Mp9@2473_d N_OUT8_Mp9@2473_g N_VDD_Mp9@2473_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2472 N_OUT9_Mp9@2472_d N_OUT8_Mp9@2472_g N_VDD_Mp9@2472_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2471 N_OUT9_Mn9@2471_d N_OUT8_Mn9@2471_g N_VSS_Mn9@2471_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2470 N_OUT9_Mn9@2470_d N_OUT8_Mn9@2470_g N_VSS_Mn9@2470_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2471 N_OUT9_Mp9@2471_d N_OUT8_Mp9@2471_g N_VDD_Mp9@2471_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2470 N_OUT9_Mp9@2470_d N_OUT8_Mp9@2470_g N_VDD_Mp9@2470_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2469 N_OUT9_Mn9@2469_d N_OUT8_Mn9@2469_g N_VSS_Mn9@2469_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2468 N_OUT9_Mn9@2468_d N_OUT8_Mn9@2468_g N_VSS_Mn9@2468_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2469 N_OUT9_Mp9@2469_d N_OUT8_Mp9@2469_g N_VDD_Mp9@2469_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2468 N_OUT9_Mp9@2468_d N_OUT8_Mp9@2468_g N_VDD_Mp9@2468_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2467 N_OUT9_Mn9@2467_d N_OUT8_Mn9@2467_g N_VSS_Mn9@2467_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2466 N_OUT9_Mn9@2466_d N_OUT8_Mn9@2466_g N_VSS_Mn9@2466_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2467 N_OUT9_Mp9@2467_d N_OUT8_Mp9@2467_g N_VDD_Mp9@2467_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2466 N_OUT9_Mp9@2466_d N_OUT8_Mp9@2466_g N_VDD_Mp9@2466_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2465 N_OUT9_Mn9@2465_d N_OUT8_Mn9@2465_g N_VSS_Mn9@2465_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2464 N_OUT9_Mn9@2464_d N_OUT8_Mn9@2464_g N_VSS_Mn9@2464_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2465 N_OUT9_Mp9@2465_d N_OUT8_Mp9@2465_g N_VDD_Mp9@2465_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2464 N_OUT9_Mp9@2464_d N_OUT8_Mp9@2464_g N_VDD_Mp9@2464_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2463 N_OUT9_Mn9@2463_d N_OUT8_Mn9@2463_g N_VSS_Mn9@2463_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2462 N_OUT9_Mn9@2462_d N_OUT8_Mn9@2462_g N_VSS_Mn9@2462_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2463 N_OUT9_Mp9@2463_d N_OUT8_Mp9@2463_g N_VDD_Mp9@2463_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2462 N_OUT9_Mp9@2462_d N_OUT8_Mp9@2462_g N_VDD_Mp9@2462_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2461 N_OUT9_Mn9@2461_d N_OUT8_Mn9@2461_g N_VSS_Mn9@2461_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2460 N_OUT9_Mn9@2460_d N_OUT8_Mn9@2460_g N_VSS_Mn9@2460_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2461 N_OUT9_Mp9@2461_d N_OUT8_Mp9@2461_g N_VDD_Mp9@2461_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2460 N_OUT9_Mp9@2460_d N_OUT8_Mp9@2460_g N_VDD_Mp9@2460_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2459 N_OUT9_Mn9@2459_d N_OUT8_Mn9@2459_g N_VSS_Mn9@2459_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2458 N_OUT9_Mn9@2458_d N_OUT8_Mn9@2458_g N_VSS_Mn9@2458_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2459 N_OUT9_Mp9@2459_d N_OUT8_Mp9@2459_g N_VDD_Mp9@2459_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2458 N_OUT9_Mp9@2458_d N_OUT8_Mp9@2458_g N_VDD_Mp9@2458_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2457 N_OUT9_Mn9@2457_d N_OUT8_Mn9@2457_g N_VSS_Mn9@2457_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2456 N_OUT9_Mn9@2456_d N_OUT8_Mn9@2456_g N_VSS_Mn9@2456_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2457 N_OUT9_Mp9@2457_d N_OUT8_Mp9@2457_g N_VDD_Mp9@2457_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2456 N_OUT9_Mp9@2456_d N_OUT8_Mp9@2456_g N_VDD_Mp9@2456_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2455 N_OUT9_Mn9@2455_d N_OUT8_Mn9@2455_g N_VSS_Mn9@2455_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2454 N_OUT9_Mn9@2454_d N_OUT8_Mn9@2454_g N_VSS_Mn9@2454_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2455 N_OUT9_Mp9@2455_d N_OUT8_Mp9@2455_g N_VDD_Mp9@2455_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2454 N_OUT9_Mp9@2454_d N_OUT8_Mp9@2454_g N_VDD_Mp9@2454_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2453 N_OUT9_Mn9@2453_d N_OUT8_Mn9@2453_g N_VSS_Mn9@2453_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2452 N_OUT9_Mn9@2452_d N_OUT8_Mn9@2452_g N_VSS_Mn9@2452_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2453 N_OUT9_Mp9@2453_d N_OUT8_Mp9@2453_g N_VDD_Mp9@2453_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2452 N_OUT9_Mp9@2452_d N_OUT8_Mp9@2452_g N_VDD_Mp9@2452_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2451 N_OUT9_Mn9@2451_d N_OUT8_Mn9@2451_g N_VSS_Mn9@2451_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2450 N_OUT9_Mn9@2450_d N_OUT8_Mn9@2450_g N_VSS_Mn9@2450_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2451 N_OUT9_Mp9@2451_d N_OUT8_Mp9@2451_g N_VDD_Mp9@2451_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2450 N_OUT9_Mp9@2450_d N_OUT8_Mp9@2450_g N_VDD_Mp9@2450_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2449 N_OUT9_Mn9@2449_d N_OUT8_Mn9@2449_g N_VSS_Mn9@2449_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2448 N_OUT9_Mn9@2448_d N_OUT8_Mn9@2448_g N_VSS_Mn9@2448_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2449 N_OUT9_Mp9@2449_d N_OUT8_Mp9@2449_g N_VDD_Mp9@2449_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2448 N_OUT9_Mp9@2448_d N_OUT8_Mp9@2448_g N_VDD_Mp9@2448_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2447 N_OUT9_Mn9@2447_d N_OUT8_Mn9@2447_g N_VSS_Mn9@2447_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2446 N_OUT9_Mn9@2446_d N_OUT8_Mn9@2446_g N_VSS_Mn9@2446_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2447 N_OUT9_Mp9@2447_d N_OUT8_Mp9@2447_g N_VDD_Mp9@2447_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2446 N_OUT9_Mp9@2446_d N_OUT8_Mp9@2446_g N_VDD_Mp9@2446_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2445 N_OUT9_Mn9@2445_d N_OUT8_Mn9@2445_g N_VSS_Mn9@2445_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2444 N_OUT9_Mn9@2444_d N_OUT8_Mn9@2444_g N_VSS_Mn9@2444_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2445 N_OUT9_Mp9@2445_d N_OUT8_Mp9@2445_g N_VDD_Mp9@2445_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2444 N_OUT9_Mp9@2444_d N_OUT8_Mp9@2444_g N_VDD_Mp9@2444_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2443 N_OUT9_Mn9@2443_d N_OUT8_Mn9@2443_g N_VSS_Mn9@2443_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2442 N_OUT9_Mn9@2442_d N_OUT8_Mn9@2442_g N_VSS_Mn9@2442_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2443 N_OUT9_Mp9@2443_d N_OUT8_Mp9@2443_g N_VDD_Mp9@2443_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2442 N_OUT9_Mp9@2442_d N_OUT8_Mp9@2442_g N_VDD_Mp9@2442_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2441 N_OUT9_Mn9@2441_d N_OUT8_Mn9@2441_g N_VSS_Mn9@2441_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2440 N_OUT9_Mn9@2440_d N_OUT8_Mn9@2440_g N_VSS_Mn9@2440_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2441 N_OUT9_Mp9@2441_d N_OUT8_Mp9@2441_g N_VDD_Mp9@2441_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2440 N_OUT9_Mp9@2440_d N_OUT8_Mp9@2440_g N_VDD_Mp9@2440_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2439 N_OUT9_Mn9@2439_d N_OUT8_Mn9@2439_g N_VSS_Mn9@2439_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2438 N_OUT9_Mn9@2438_d N_OUT8_Mn9@2438_g N_VSS_Mn9@2438_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2439 N_OUT9_Mp9@2439_d N_OUT8_Mp9@2439_g N_VDD_Mp9@2439_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2438 N_OUT9_Mp9@2438_d N_OUT8_Mp9@2438_g N_VDD_Mp9@2438_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2437 N_OUT9_Mn9@2437_d N_OUT8_Mn9@2437_g N_VSS_Mn9@2437_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2436 N_OUT9_Mn9@2436_d N_OUT8_Mn9@2436_g N_VSS_Mn9@2436_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2437 N_OUT9_Mp9@2437_d N_OUT8_Mp9@2437_g N_VDD_Mp9@2437_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2436 N_OUT9_Mp9@2436_d N_OUT8_Mp9@2436_g N_VDD_Mp9@2436_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2435 N_OUT9_Mn9@2435_d N_OUT8_Mn9@2435_g N_VSS_Mn9@2435_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2434 N_OUT9_Mn9@2434_d N_OUT8_Mn9@2434_g N_VSS_Mn9@2434_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2435 N_OUT9_Mp9@2435_d N_OUT8_Mp9@2435_g N_VDD_Mp9@2435_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2434 N_OUT9_Mp9@2434_d N_OUT8_Mp9@2434_g N_VDD_Mp9@2434_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2433 N_OUT9_Mn9@2433_d N_OUT8_Mn9@2433_g N_VSS_Mn9@2433_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2432 N_OUT9_Mn9@2432_d N_OUT8_Mn9@2432_g N_VSS_Mn9@2432_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2433 N_OUT9_Mp9@2433_d N_OUT8_Mp9@2433_g N_VDD_Mp9@2433_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2432 N_OUT9_Mp9@2432_d N_OUT8_Mp9@2432_g N_VDD_Mp9@2432_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2431 N_OUT9_Mn9@2431_d N_OUT8_Mn9@2431_g N_VSS_Mn9@2431_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2430 N_OUT9_Mn9@2430_d N_OUT8_Mn9@2430_g N_VSS_Mn9@2430_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2431 N_OUT9_Mp9@2431_d N_OUT8_Mp9@2431_g N_VDD_Mp9@2431_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2430 N_OUT9_Mp9@2430_d N_OUT8_Mp9@2430_g N_VDD_Mp9@2430_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2429 N_OUT9_Mn9@2429_d N_OUT8_Mn9@2429_g N_VSS_Mn9@2429_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2428 N_OUT9_Mn9@2428_d N_OUT8_Mn9@2428_g N_VSS_Mn9@2428_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2429 N_OUT9_Mp9@2429_d N_OUT8_Mp9@2429_g N_VDD_Mp9@2429_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2428 N_OUT9_Mp9@2428_d N_OUT8_Mp9@2428_g N_VDD_Mp9@2428_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2427 N_OUT9_Mn9@2427_d N_OUT8_Mn9@2427_g N_VSS_Mn9@2427_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2426 N_OUT9_Mn9@2426_d N_OUT8_Mn9@2426_g N_VSS_Mn9@2426_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2427 N_OUT9_Mp9@2427_d N_OUT8_Mp9@2427_g N_VDD_Mp9@2427_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2426 N_OUT9_Mp9@2426_d N_OUT8_Mp9@2426_g N_VDD_Mp9@2426_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2425 N_OUT9_Mn9@2425_d N_OUT8_Mn9@2425_g N_VSS_Mn9@2425_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2424 N_OUT9_Mn9@2424_d N_OUT8_Mn9@2424_g N_VSS_Mn9@2424_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2425 N_OUT9_Mp9@2425_d N_OUT8_Mp9@2425_g N_VDD_Mp9@2425_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2424 N_OUT9_Mp9@2424_d N_OUT8_Mp9@2424_g N_VDD_Mp9@2424_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2423 N_OUT9_Mn9@2423_d N_OUT8_Mn9@2423_g N_VSS_Mn9@2423_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2422 N_OUT9_Mn9@2422_d N_OUT8_Mn9@2422_g N_VSS_Mn9@2422_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2423 N_OUT9_Mp9@2423_d N_OUT8_Mp9@2423_g N_VDD_Mp9@2423_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2422 N_OUT9_Mp9@2422_d N_OUT8_Mp9@2422_g N_VDD_Mp9@2422_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2421 N_OUT9_Mn9@2421_d N_OUT8_Mn9@2421_g N_VSS_Mn9@2421_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2420 N_OUT9_Mn9@2420_d N_OUT8_Mn9@2420_g N_VSS_Mn9@2420_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2421 N_OUT9_Mp9@2421_d N_OUT8_Mp9@2421_g N_VDD_Mp9@2421_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2420 N_OUT9_Mp9@2420_d N_OUT8_Mp9@2420_g N_VDD_Mp9@2420_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2419 N_OUT9_Mn9@2419_d N_OUT8_Mn9@2419_g N_VSS_Mn9@2419_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2418 N_OUT9_Mn9@2418_d N_OUT8_Mn9@2418_g N_VSS_Mn9@2418_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2419 N_OUT9_Mp9@2419_d N_OUT8_Mp9@2419_g N_VDD_Mp9@2419_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2418 N_OUT9_Mp9@2418_d N_OUT8_Mp9@2418_g N_VDD_Mp9@2418_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2417 N_OUT9_Mn9@2417_d N_OUT8_Mn9@2417_g N_VSS_Mn9@2417_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2416 N_OUT9_Mn9@2416_d N_OUT8_Mn9@2416_g N_VSS_Mn9@2416_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2417 N_OUT9_Mp9@2417_d N_OUT8_Mp9@2417_g N_VDD_Mp9@2417_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2416 N_OUT9_Mp9@2416_d N_OUT8_Mp9@2416_g N_VDD_Mp9@2416_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2415 N_OUT9_Mn9@2415_d N_OUT8_Mn9@2415_g N_VSS_Mn9@2415_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2414 N_OUT9_Mn9@2414_d N_OUT8_Mn9@2414_g N_VSS_Mn9@2414_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2415 N_OUT9_Mp9@2415_d N_OUT8_Mp9@2415_g N_VDD_Mp9@2415_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2414 N_OUT9_Mp9@2414_d N_OUT8_Mp9@2414_g N_VDD_Mp9@2414_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2413 N_OUT9_Mn9@2413_d N_OUT8_Mn9@2413_g N_VSS_Mn9@2413_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2412 N_OUT9_Mn9@2412_d N_OUT8_Mn9@2412_g N_VSS_Mn9@2412_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2413 N_OUT9_Mp9@2413_d N_OUT8_Mp9@2413_g N_VDD_Mp9@2413_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2412 N_OUT9_Mp9@2412_d N_OUT8_Mp9@2412_g N_VDD_Mp9@2412_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2411 N_OUT9_Mn9@2411_d N_OUT8_Mn9@2411_g N_VSS_Mn9@2411_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2410 N_OUT9_Mn9@2410_d N_OUT8_Mn9@2410_g N_VSS_Mn9@2410_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2411 N_OUT9_Mp9@2411_d N_OUT8_Mp9@2411_g N_VDD_Mp9@2411_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2410 N_OUT9_Mp9@2410_d N_OUT8_Mp9@2410_g N_VDD_Mp9@2410_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2409 N_OUT9_Mn9@2409_d N_OUT8_Mn9@2409_g N_VSS_Mn9@2409_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2408 N_OUT9_Mn9@2408_d N_OUT8_Mn9@2408_g N_VSS_Mn9@2408_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2409 N_OUT9_Mp9@2409_d N_OUT8_Mp9@2409_g N_VDD_Mp9@2409_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2408 N_OUT9_Mp9@2408_d N_OUT8_Mp9@2408_g N_VDD_Mp9@2408_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2407 N_OUT9_Mn9@2407_d N_OUT8_Mn9@2407_g N_VSS_Mn9@2407_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2406 N_OUT9_Mn9@2406_d N_OUT8_Mn9@2406_g N_VSS_Mn9@2406_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2407 N_OUT9_Mp9@2407_d N_OUT8_Mp9@2407_g N_VDD_Mp9@2407_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2406 N_OUT9_Mp9@2406_d N_OUT8_Mp9@2406_g N_VDD_Mp9@2406_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2405 N_OUT9_Mn9@2405_d N_OUT8_Mn9@2405_g N_VSS_Mn9@2405_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2404 N_OUT9_Mn9@2404_d N_OUT8_Mn9@2404_g N_VSS_Mn9@2404_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2405 N_OUT9_Mp9@2405_d N_OUT8_Mp9@2405_g N_VDD_Mp9@2405_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2404 N_OUT9_Mp9@2404_d N_OUT8_Mp9@2404_g N_VDD_Mp9@2404_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2403 N_OUT9_Mn9@2403_d N_OUT8_Mn9@2403_g N_VSS_Mn9@2403_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2402 N_OUT9_Mn9@2402_d N_OUT8_Mn9@2402_g N_VSS_Mn9@2402_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2403 N_OUT9_Mp9@2403_d N_OUT8_Mp9@2403_g N_VDD_Mp9@2403_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2402 N_OUT9_Mp9@2402_d N_OUT8_Mp9@2402_g N_VDD_Mp9@2402_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2401 N_OUT9_Mn9@2401_d N_OUT8_Mn9@2401_g N_VSS_Mn9@2401_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2400 N_OUT9_Mn9@2400_d N_OUT8_Mn9@2400_g N_VSS_Mn9@2400_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2401 N_OUT9_Mp9@2401_d N_OUT8_Mp9@2401_g N_VDD_Mp9@2401_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2400 N_OUT9_Mp9@2400_d N_OUT8_Mp9@2400_g N_VDD_Mp9@2400_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2399 N_OUT9_Mn9@2399_d N_OUT8_Mn9@2399_g N_VSS_Mn9@2399_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2398 N_OUT9_Mn9@2398_d N_OUT8_Mn9@2398_g N_VSS_Mn9@2398_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2399 N_OUT9_Mp9@2399_d N_OUT8_Mp9@2399_g N_VDD_Mp9@2399_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2398 N_OUT9_Mp9@2398_d N_OUT8_Mp9@2398_g N_VDD_Mp9@2398_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2397 N_OUT9_Mn9@2397_d N_OUT8_Mn9@2397_g N_VSS_Mn9@2397_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2396 N_OUT9_Mn9@2396_d N_OUT8_Mn9@2396_g N_VSS_Mn9@2396_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2397 N_OUT9_Mp9@2397_d N_OUT8_Mp9@2397_g N_VDD_Mp9@2397_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2396 N_OUT9_Mp9@2396_d N_OUT8_Mp9@2396_g N_VDD_Mp9@2396_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2395 N_OUT9_Mn9@2395_d N_OUT8_Mn9@2395_g N_VSS_Mn9@2395_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2394 N_OUT9_Mn9@2394_d N_OUT8_Mn9@2394_g N_VSS_Mn9@2394_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2395 N_OUT9_Mp9@2395_d N_OUT8_Mp9@2395_g N_VDD_Mp9@2395_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2394 N_OUT9_Mp9@2394_d N_OUT8_Mp9@2394_g N_VDD_Mp9@2394_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2393 N_OUT9_Mn9@2393_d N_OUT8_Mn9@2393_g N_VSS_Mn9@2393_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2392 N_OUT9_Mn9@2392_d N_OUT8_Mn9@2392_g N_VSS_Mn9@2392_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2393 N_OUT9_Mp9@2393_d N_OUT8_Mp9@2393_g N_VDD_Mp9@2393_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2392 N_OUT9_Mp9@2392_d N_OUT8_Mp9@2392_g N_VDD_Mp9@2392_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2391 N_OUT9_Mn9@2391_d N_OUT8_Mn9@2391_g N_VSS_Mn9@2391_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2390 N_OUT9_Mn9@2390_d N_OUT8_Mn9@2390_g N_VSS_Mn9@2390_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2391 N_OUT9_Mp9@2391_d N_OUT8_Mp9@2391_g N_VDD_Mp9@2391_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2390 N_OUT9_Mp9@2390_d N_OUT8_Mp9@2390_g N_VDD_Mp9@2390_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2389 N_OUT9_Mn9@2389_d N_OUT8_Mn9@2389_g N_VSS_Mn9@2389_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2388 N_OUT9_Mn9@2388_d N_OUT8_Mn9@2388_g N_VSS_Mn9@2388_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2389 N_OUT9_Mp9@2389_d N_OUT8_Mp9@2389_g N_VDD_Mp9@2389_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2388 N_OUT9_Mp9@2388_d N_OUT8_Mp9@2388_g N_VDD_Mp9@2388_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2387 N_OUT9_Mn9@2387_d N_OUT8_Mn9@2387_g N_VSS_Mn9@2387_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2386 N_OUT9_Mn9@2386_d N_OUT8_Mn9@2386_g N_VSS_Mn9@2386_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2387 N_OUT9_Mp9@2387_d N_OUT8_Mp9@2387_g N_VDD_Mp9@2387_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2386 N_OUT9_Mp9@2386_d N_OUT8_Mp9@2386_g N_VDD_Mp9@2386_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2385 N_OUT9_Mn9@2385_d N_OUT8_Mn9@2385_g N_VSS_Mn9@2385_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2384 N_OUT9_Mn9@2384_d N_OUT8_Mn9@2384_g N_VSS_Mn9@2384_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2385 N_OUT9_Mp9@2385_d N_OUT8_Mp9@2385_g N_VDD_Mp9@2385_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2384 N_OUT9_Mp9@2384_d N_OUT8_Mp9@2384_g N_VDD_Mp9@2384_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2383 N_OUT9_Mn9@2383_d N_OUT8_Mn9@2383_g N_VSS_Mn9@2383_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2382 N_OUT9_Mn9@2382_d N_OUT8_Mn9@2382_g N_VSS_Mn9@2382_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2383 N_OUT9_Mp9@2383_d N_OUT8_Mp9@2383_g N_VDD_Mp9@2383_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2382 N_OUT9_Mp9@2382_d N_OUT8_Mp9@2382_g N_VDD_Mp9@2382_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2381 N_OUT9_Mn9@2381_d N_OUT8_Mn9@2381_g N_VSS_Mn9@2381_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2380 N_OUT9_Mn9@2380_d N_OUT8_Mn9@2380_g N_VSS_Mn9@2380_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2381 N_OUT9_Mp9@2381_d N_OUT8_Mp9@2381_g N_VDD_Mp9@2381_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2380 N_OUT9_Mp9@2380_d N_OUT8_Mp9@2380_g N_VDD_Mp9@2380_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2379 N_OUT9_Mn9@2379_d N_OUT8_Mn9@2379_g N_VSS_Mn9@2379_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2378 N_OUT9_Mn9@2378_d N_OUT8_Mn9@2378_g N_VSS_Mn9@2378_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2379 N_OUT9_Mp9@2379_d N_OUT8_Mp9@2379_g N_VDD_Mp9@2379_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2378 N_OUT9_Mp9@2378_d N_OUT8_Mp9@2378_g N_VDD_Mp9@2378_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2377 N_OUT9_Mn9@2377_d N_OUT8_Mn9@2377_g N_VSS_Mn9@2377_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2376 N_OUT9_Mn9@2376_d N_OUT8_Mn9@2376_g N_VSS_Mn9@2376_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2377 N_OUT9_Mp9@2377_d N_OUT8_Mp9@2377_g N_VDD_Mp9@2377_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2376 N_OUT9_Mp9@2376_d N_OUT8_Mp9@2376_g N_VDD_Mp9@2376_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2375 N_OUT9_Mn9@2375_d N_OUT8_Mn9@2375_g N_VSS_Mn9@2375_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2374 N_OUT9_Mn9@2374_d N_OUT8_Mn9@2374_g N_VSS_Mn9@2374_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2375 N_OUT9_Mp9@2375_d N_OUT8_Mp9@2375_g N_VDD_Mp9@2375_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2374 N_OUT9_Mp9@2374_d N_OUT8_Mp9@2374_g N_VDD_Mp9@2374_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2373 N_OUT9_Mn9@2373_d N_OUT8_Mn9@2373_g N_VSS_Mn9@2373_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2372 N_OUT9_Mn9@2372_d N_OUT8_Mn9@2372_g N_VSS_Mn9@2372_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2373 N_OUT9_Mp9@2373_d N_OUT8_Mp9@2373_g N_VDD_Mp9@2373_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2372 N_OUT9_Mp9@2372_d N_OUT8_Mp9@2372_g N_VDD_Mp9@2372_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2371 N_OUT9_Mn9@2371_d N_OUT8_Mn9@2371_g N_VSS_Mn9@2371_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2370 N_OUT9_Mn9@2370_d N_OUT8_Mn9@2370_g N_VSS_Mn9@2370_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2371 N_OUT9_Mp9@2371_d N_OUT8_Mp9@2371_g N_VDD_Mp9@2371_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2370 N_OUT9_Mp9@2370_d N_OUT8_Mp9@2370_g N_VDD_Mp9@2370_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2369 N_OUT9_Mn9@2369_d N_OUT8_Mn9@2369_g N_VSS_Mn9@2369_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2368 N_OUT9_Mn9@2368_d N_OUT8_Mn9@2368_g N_VSS_Mn9@2368_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2369 N_OUT9_Mp9@2369_d N_OUT8_Mp9@2369_g N_VDD_Mp9@2369_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2368 N_OUT9_Mp9@2368_d N_OUT8_Mp9@2368_g N_VDD_Mp9@2368_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2367 N_OUT9_Mn9@2367_d N_OUT8_Mn9@2367_g N_VSS_Mn9@2367_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2366 N_OUT9_Mn9@2366_d N_OUT8_Mn9@2366_g N_VSS_Mn9@2366_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2367 N_OUT9_Mp9@2367_d N_OUT8_Mp9@2367_g N_VDD_Mp9@2367_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2366 N_OUT9_Mp9@2366_d N_OUT8_Mp9@2366_g N_VDD_Mp9@2366_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2365 N_OUT9_Mn9@2365_d N_OUT8_Mn9@2365_g N_VSS_Mn9@2365_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2364 N_OUT9_Mn9@2364_d N_OUT8_Mn9@2364_g N_VSS_Mn9@2364_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2365 N_OUT9_Mp9@2365_d N_OUT8_Mp9@2365_g N_VDD_Mp9@2365_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2364 N_OUT9_Mp9@2364_d N_OUT8_Mp9@2364_g N_VDD_Mp9@2364_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2363 N_OUT9_Mn9@2363_d N_OUT8_Mn9@2363_g N_VSS_Mn9@2363_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2362 N_OUT9_Mn9@2362_d N_OUT8_Mn9@2362_g N_VSS_Mn9@2362_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2363 N_OUT9_Mp9@2363_d N_OUT8_Mp9@2363_g N_VDD_Mp9@2363_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2362 N_OUT9_Mp9@2362_d N_OUT8_Mp9@2362_g N_VDD_Mp9@2362_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2361 N_OUT9_Mn9@2361_d N_OUT8_Mn9@2361_g N_VSS_Mn9@2361_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2360 N_OUT9_Mn9@2360_d N_OUT8_Mn9@2360_g N_VSS_Mn9@2360_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2361 N_OUT9_Mp9@2361_d N_OUT8_Mp9@2361_g N_VDD_Mp9@2361_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2360 N_OUT9_Mp9@2360_d N_OUT8_Mp9@2360_g N_VDD_Mp9@2360_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2359 N_OUT9_Mn9@2359_d N_OUT8_Mn9@2359_g N_VSS_Mn9@2359_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2358 N_OUT9_Mn9@2358_d N_OUT8_Mn9@2358_g N_VSS_Mn9@2358_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2359 N_OUT9_Mp9@2359_d N_OUT8_Mp9@2359_g N_VDD_Mp9@2359_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2358 N_OUT9_Mp9@2358_d N_OUT8_Mp9@2358_g N_VDD_Mp9@2358_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2357 N_OUT9_Mn9@2357_d N_OUT8_Mn9@2357_g N_VSS_Mn9@2357_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2356 N_OUT9_Mn9@2356_d N_OUT8_Mn9@2356_g N_VSS_Mn9@2356_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2357 N_OUT9_Mp9@2357_d N_OUT8_Mp9@2357_g N_VDD_Mp9@2357_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2356 N_OUT9_Mp9@2356_d N_OUT8_Mp9@2356_g N_VDD_Mp9@2356_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2355 N_OUT9_Mn9@2355_d N_OUT8_Mn9@2355_g N_VSS_Mn9@2355_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2354 N_OUT9_Mn9@2354_d N_OUT8_Mn9@2354_g N_VSS_Mn9@2354_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2355 N_OUT9_Mp9@2355_d N_OUT8_Mp9@2355_g N_VDD_Mp9@2355_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2354 N_OUT9_Mp9@2354_d N_OUT8_Mp9@2354_g N_VDD_Mp9@2354_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2353 N_OUT9_Mn9@2353_d N_OUT8_Mn9@2353_g N_VSS_Mn9@2353_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2352 N_OUT9_Mn9@2352_d N_OUT8_Mn9@2352_g N_VSS_Mn9@2352_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2353 N_OUT9_Mp9@2353_d N_OUT8_Mp9@2353_g N_VDD_Mp9@2353_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2352 N_OUT9_Mp9@2352_d N_OUT8_Mp9@2352_g N_VDD_Mp9@2352_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2351 N_OUT9_Mn9@2351_d N_OUT8_Mn9@2351_g N_VSS_Mn9@2351_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2350 N_OUT9_Mn9@2350_d N_OUT8_Mn9@2350_g N_VSS_Mn9@2350_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2351 N_OUT9_Mp9@2351_d N_OUT8_Mp9@2351_g N_VDD_Mp9@2351_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2350 N_OUT9_Mp9@2350_d N_OUT8_Mp9@2350_g N_VDD_Mp9@2350_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2349 N_OUT9_Mn9@2349_d N_OUT8_Mn9@2349_g N_VSS_Mn9@2349_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2348 N_OUT9_Mn9@2348_d N_OUT8_Mn9@2348_g N_VSS_Mn9@2348_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2349 N_OUT9_Mp9@2349_d N_OUT8_Mp9@2349_g N_VDD_Mp9@2349_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2348 N_OUT9_Mp9@2348_d N_OUT8_Mp9@2348_g N_VDD_Mp9@2348_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2347 N_OUT9_Mn9@2347_d N_OUT8_Mn9@2347_g N_VSS_Mn9@2347_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2346 N_OUT9_Mn9@2346_d N_OUT8_Mn9@2346_g N_VSS_Mn9@2346_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2347 N_OUT9_Mp9@2347_d N_OUT8_Mp9@2347_g N_VDD_Mp9@2347_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2346 N_OUT9_Mp9@2346_d N_OUT8_Mp9@2346_g N_VDD_Mp9@2346_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2345 N_OUT9_Mn9@2345_d N_OUT8_Mn9@2345_g N_VSS_Mn9@2345_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2344 N_OUT9_Mn9@2344_d N_OUT8_Mn9@2344_g N_VSS_Mn9@2344_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2345 N_OUT9_Mp9@2345_d N_OUT8_Mp9@2345_g N_VDD_Mp9@2345_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2344 N_OUT9_Mp9@2344_d N_OUT8_Mp9@2344_g N_VDD_Mp9@2344_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2343 N_OUT9_Mn9@2343_d N_OUT8_Mn9@2343_g N_VSS_Mn9@2343_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2342 N_OUT9_Mn9@2342_d N_OUT8_Mn9@2342_g N_VSS_Mn9@2342_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2343 N_OUT9_Mp9@2343_d N_OUT8_Mp9@2343_g N_VDD_Mp9@2343_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2342 N_OUT9_Mp9@2342_d N_OUT8_Mp9@2342_g N_VDD_Mp9@2342_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2341 N_OUT9_Mn9@2341_d N_OUT8_Mn9@2341_g N_VSS_Mn9@2341_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2340 N_OUT9_Mn9@2340_d N_OUT8_Mn9@2340_g N_VSS_Mn9@2340_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2341 N_OUT9_Mp9@2341_d N_OUT8_Mp9@2341_g N_VDD_Mp9@2341_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2340 N_OUT9_Mp9@2340_d N_OUT8_Mp9@2340_g N_VDD_Mp9@2340_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2339 N_OUT9_Mn9@2339_d N_OUT8_Mn9@2339_g N_VSS_Mn9@2339_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2338 N_OUT9_Mn9@2338_d N_OUT8_Mn9@2338_g N_VSS_Mn9@2338_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2339 N_OUT9_Mp9@2339_d N_OUT8_Mp9@2339_g N_VDD_Mp9@2339_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2338 N_OUT9_Mp9@2338_d N_OUT8_Mp9@2338_g N_VDD_Mp9@2338_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2337 N_OUT9_Mn9@2337_d N_OUT8_Mn9@2337_g N_VSS_Mn9@2337_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2336 N_OUT9_Mn9@2336_d N_OUT8_Mn9@2336_g N_VSS_Mn9@2336_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2337 N_OUT9_Mp9@2337_d N_OUT8_Mp9@2337_g N_VDD_Mp9@2337_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2336 N_OUT9_Mp9@2336_d N_OUT8_Mp9@2336_g N_VDD_Mp9@2336_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2335 N_OUT9_Mn9@2335_d N_OUT8_Mn9@2335_g N_VSS_Mn9@2335_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2334 N_OUT9_Mn9@2334_d N_OUT8_Mn9@2334_g N_VSS_Mn9@2334_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2335 N_OUT9_Mp9@2335_d N_OUT8_Mp9@2335_g N_VDD_Mp9@2335_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2334 N_OUT9_Mp9@2334_d N_OUT8_Mp9@2334_g N_VDD_Mp9@2334_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2333 N_OUT9_Mn9@2333_d N_OUT8_Mn9@2333_g N_VSS_Mn9@2333_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2332 N_OUT9_Mn9@2332_d N_OUT8_Mn9@2332_g N_VSS_Mn9@2332_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2333 N_OUT9_Mp9@2333_d N_OUT8_Mp9@2333_g N_VDD_Mp9@2333_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2332 N_OUT9_Mp9@2332_d N_OUT8_Mp9@2332_g N_VDD_Mp9@2332_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2331 N_OUT9_Mn9@2331_d N_OUT8_Mn9@2331_g N_VSS_Mn9@2331_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2330 N_OUT9_Mn9@2330_d N_OUT8_Mn9@2330_g N_VSS_Mn9@2330_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2331 N_OUT9_Mp9@2331_d N_OUT8_Mp9@2331_g N_VDD_Mp9@2331_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2330 N_OUT9_Mp9@2330_d N_OUT8_Mp9@2330_g N_VDD_Mp9@2330_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2329 N_OUT9_Mn9@2329_d N_OUT8_Mn9@2329_g N_VSS_Mn9@2329_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2328 N_OUT9_Mn9@2328_d N_OUT8_Mn9@2328_g N_VSS_Mn9@2328_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2329 N_OUT9_Mp9@2329_d N_OUT8_Mp9@2329_g N_VDD_Mp9@2329_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2328 N_OUT9_Mp9@2328_d N_OUT8_Mp9@2328_g N_VDD_Mp9@2328_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2327 N_OUT9_Mn9@2327_d N_OUT8_Mn9@2327_g N_VSS_Mn9@2327_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2326 N_OUT9_Mn9@2326_d N_OUT8_Mn9@2326_g N_VSS_Mn9@2326_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2327 N_OUT9_Mp9@2327_d N_OUT8_Mp9@2327_g N_VDD_Mp9@2327_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2326 N_OUT9_Mp9@2326_d N_OUT8_Mp9@2326_g N_VDD_Mp9@2326_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2325 N_OUT9_Mn9@2325_d N_OUT8_Mn9@2325_g N_VSS_Mn9@2325_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2324 N_OUT9_Mn9@2324_d N_OUT8_Mn9@2324_g N_VSS_Mn9@2324_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2325 N_OUT9_Mp9@2325_d N_OUT8_Mp9@2325_g N_VDD_Mp9@2325_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2324 N_OUT9_Mp9@2324_d N_OUT8_Mp9@2324_g N_VDD_Mp9@2324_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2323 N_OUT9_Mn9@2323_d N_OUT8_Mn9@2323_g N_VSS_Mn9@2323_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2322 N_OUT9_Mn9@2322_d N_OUT8_Mn9@2322_g N_VSS_Mn9@2322_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2323 N_OUT9_Mp9@2323_d N_OUT8_Mp9@2323_g N_VDD_Mp9@2323_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2322 N_OUT9_Mp9@2322_d N_OUT8_Mp9@2322_g N_VDD_Mp9@2322_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2321 N_OUT9_Mn9@2321_d N_OUT8_Mn9@2321_g N_VSS_Mn9@2321_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2320 N_OUT9_Mn9@2320_d N_OUT8_Mn9@2320_g N_VSS_Mn9@2320_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2321 N_OUT9_Mp9@2321_d N_OUT8_Mp9@2321_g N_VDD_Mp9@2321_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2320 N_OUT9_Mp9@2320_d N_OUT8_Mp9@2320_g N_VDD_Mp9@2320_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2319 N_OUT9_Mn9@2319_d N_OUT8_Mn9@2319_g N_VSS_Mn9@2319_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2318 N_OUT9_Mn9@2318_d N_OUT8_Mn9@2318_g N_VSS_Mn9@2318_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2319 N_OUT9_Mp9@2319_d N_OUT8_Mp9@2319_g N_VDD_Mp9@2319_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2318 N_OUT9_Mp9@2318_d N_OUT8_Mp9@2318_g N_VDD_Mp9@2318_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2317 N_OUT9_Mn9@2317_d N_OUT8_Mn9@2317_g N_VSS_Mn9@2317_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2316 N_OUT9_Mn9@2316_d N_OUT8_Mn9@2316_g N_VSS_Mn9@2316_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2317 N_OUT9_Mp9@2317_d N_OUT8_Mp9@2317_g N_VDD_Mp9@2317_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2316 N_OUT9_Mp9@2316_d N_OUT8_Mp9@2316_g N_VDD_Mp9@2316_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2315 N_OUT9_Mn9@2315_d N_OUT8_Mn9@2315_g N_VSS_Mn9@2315_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2314 N_OUT9_Mn9@2314_d N_OUT8_Mn9@2314_g N_VSS_Mn9@2314_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2315 N_OUT9_Mp9@2315_d N_OUT8_Mp9@2315_g N_VDD_Mp9@2315_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2314 N_OUT9_Mp9@2314_d N_OUT8_Mp9@2314_g N_VDD_Mp9@2314_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2313 N_OUT9_Mn9@2313_d N_OUT8_Mn9@2313_g N_VSS_Mn9@2313_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2312 N_OUT9_Mn9@2312_d N_OUT8_Mn9@2312_g N_VSS_Mn9@2312_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2313 N_OUT9_Mp9@2313_d N_OUT8_Mp9@2313_g N_VDD_Mp9@2313_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2312 N_OUT9_Mp9@2312_d N_OUT8_Mp9@2312_g N_VDD_Mp9@2312_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2311 N_OUT9_Mn9@2311_d N_OUT8_Mn9@2311_g N_VSS_Mn9@2311_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2310 N_OUT9_Mn9@2310_d N_OUT8_Mn9@2310_g N_VSS_Mn9@2310_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2311 N_OUT9_Mp9@2311_d N_OUT8_Mp9@2311_g N_VDD_Mp9@2311_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2310 N_OUT9_Mp9@2310_d N_OUT8_Mp9@2310_g N_VDD_Mp9@2310_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2309 N_OUT9_Mn9@2309_d N_OUT8_Mn9@2309_g N_VSS_Mn9@2309_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2308 N_OUT9_Mn9@2308_d N_OUT8_Mn9@2308_g N_VSS_Mn9@2308_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2309 N_OUT9_Mp9@2309_d N_OUT8_Mp9@2309_g N_VDD_Mp9@2309_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2308 N_OUT9_Mp9@2308_d N_OUT8_Mp9@2308_g N_VDD_Mp9@2308_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2307 N_OUT9_Mn9@2307_d N_OUT8_Mn9@2307_g N_VSS_Mn9@2307_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2306 N_OUT9_Mn9@2306_d N_OUT8_Mn9@2306_g N_VSS_Mn9@2306_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2307 N_OUT9_Mp9@2307_d N_OUT8_Mp9@2307_g N_VDD_Mp9@2307_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2306 N_OUT9_Mp9@2306_d N_OUT8_Mp9@2306_g N_VDD_Mp9@2306_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2305 N_OUT9_Mn9@2305_d N_OUT8_Mn9@2305_g N_VSS_Mn9@2305_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2304 N_OUT9_Mn9@2304_d N_OUT8_Mn9@2304_g N_VSS_Mn9@2304_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2305 N_OUT9_Mp9@2305_d N_OUT8_Mp9@2305_g N_VDD_Mp9@2305_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2304 N_OUT9_Mp9@2304_d N_OUT8_Mp9@2304_g N_VDD_Mp9@2304_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2303 N_OUT9_Mn9@2303_d N_OUT8_Mn9@2303_g N_VSS_Mn9@2303_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2302 N_OUT9_Mn9@2302_d N_OUT8_Mn9@2302_g N_VSS_Mn9@2302_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2303 N_OUT9_Mp9@2303_d N_OUT8_Mp9@2303_g N_VDD_Mp9@2303_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2302 N_OUT9_Mp9@2302_d N_OUT8_Mp9@2302_g N_VDD_Mp9@2302_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2301 N_OUT9_Mn9@2301_d N_OUT8_Mn9@2301_g N_VSS_Mn9@2301_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2300 N_OUT9_Mn9@2300_d N_OUT8_Mn9@2300_g N_VSS_Mn9@2300_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2301 N_OUT9_Mp9@2301_d N_OUT8_Mp9@2301_g N_VDD_Mp9@2301_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2300 N_OUT9_Mp9@2300_d N_OUT8_Mp9@2300_g N_VDD_Mp9@2300_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2299 N_OUT9_Mn9@2299_d N_OUT8_Mn9@2299_g N_VSS_Mn9@2299_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2298 N_OUT9_Mn9@2298_d N_OUT8_Mn9@2298_g N_VSS_Mn9@2298_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2299 N_OUT9_Mp9@2299_d N_OUT8_Mp9@2299_g N_VDD_Mp9@2299_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2298 N_OUT9_Mp9@2298_d N_OUT8_Mp9@2298_g N_VDD_Mp9@2298_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2297 N_OUT9_Mn9@2297_d N_OUT8_Mn9@2297_g N_VSS_Mn9@2297_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2296 N_OUT9_Mn9@2296_d N_OUT8_Mn9@2296_g N_VSS_Mn9@2296_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2297 N_OUT9_Mp9@2297_d N_OUT8_Mp9@2297_g N_VDD_Mp9@2297_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2296 N_OUT9_Mp9@2296_d N_OUT8_Mp9@2296_g N_VDD_Mp9@2296_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2295 N_OUT9_Mn9@2295_d N_OUT8_Mn9@2295_g N_VSS_Mn9@2295_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2294 N_OUT9_Mn9@2294_d N_OUT8_Mn9@2294_g N_VSS_Mn9@2294_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2295 N_OUT9_Mp9@2295_d N_OUT8_Mp9@2295_g N_VDD_Mp9@2295_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2294 N_OUT9_Mp9@2294_d N_OUT8_Mp9@2294_g N_VDD_Mp9@2294_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2293 N_OUT9_Mn9@2293_d N_OUT8_Mn9@2293_g N_VSS_Mn9@2293_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2292 N_OUT9_Mn9@2292_d N_OUT8_Mn9@2292_g N_VSS_Mn9@2292_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2293 N_OUT9_Mp9@2293_d N_OUT8_Mp9@2293_g N_VDD_Mp9@2293_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2292 N_OUT9_Mp9@2292_d N_OUT8_Mp9@2292_g N_VDD_Mp9@2292_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2291 N_OUT9_Mn9@2291_d N_OUT8_Mn9@2291_g N_VSS_Mn9@2291_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2290 N_OUT9_Mn9@2290_d N_OUT8_Mn9@2290_g N_VSS_Mn9@2290_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2291 N_OUT9_Mp9@2291_d N_OUT8_Mp9@2291_g N_VDD_Mp9@2291_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2290 N_OUT9_Mp9@2290_d N_OUT8_Mp9@2290_g N_VDD_Mp9@2290_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2289 N_OUT9_Mn9@2289_d N_OUT8_Mn9@2289_g N_VSS_Mn9@2289_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2288 N_OUT9_Mn9@2288_d N_OUT8_Mn9@2288_g N_VSS_Mn9@2288_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2289 N_OUT9_Mp9@2289_d N_OUT8_Mp9@2289_g N_VDD_Mp9@2289_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2288 N_OUT9_Mp9@2288_d N_OUT8_Mp9@2288_g N_VDD_Mp9@2288_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2287 N_OUT9_Mn9@2287_d N_OUT8_Mn9@2287_g N_VSS_Mn9@2287_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2286 N_OUT9_Mn9@2286_d N_OUT8_Mn9@2286_g N_VSS_Mn9@2286_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2287 N_OUT9_Mp9@2287_d N_OUT8_Mp9@2287_g N_VDD_Mp9@2287_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2286 N_OUT9_Mp9@2286_d N_OUT8_Mp9@2286_g N_VDD_Mp9@2286_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2285 N_OUT9_Mn9@2285_d N_OUT8_Mn9@2285_g N_VSS_Mn9@2285_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2284 N_OUT9_Mn9@2284_d N_OUT8_Mn9@2284_g N_VSS_Mn9@2284_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2285 N_OUT9_Mp9@2285_d N_OUT8_Mp9@2285_g N_VDD_Mp9@2285_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2284 N_OUT9_Mp9@2284_d N_OUT8_Mp9@2284_g N_VDD_Mp9@2284_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2283 N_OUT9_Mn9@2283_d N_OUT8_Mn9@2283_g N_VSS_Mn9@2283_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2282 N_OUT9_Mn9@2282_d N_OUT8_Mn9@2282_g N_VSS_Mn9@2282_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2283 N_OUT9_Mp9@2283_d N_OUT8_Mp9@2283_g N_VDD_Mp9@2283_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2282 N_OUT9_Mp9@2282_d N_OUT8_Mp9@2282_g N_VDD_Mp9@2282_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2281 N_OUT9_Mn9@2281_d N_OUT8_Mn9@2281_g N_VSS_Mn9@2281_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2280 N_OUT9_Mn9@2280_d N_OUT8_Mn9@2280_g N_VSS_Mn9@2280_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2281 N_OUT9_Mp9@2281_d N_OUT8_Mp9@2281_g N_VDD_Mp9@2281_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2280 N_OUT9_Mp9@2280_d N_OUT8_Mp9@2280_g N_VDD_Mp9@2280_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2279 N_OUT9_Mn9@2279_d N_OUT8_Mn9@2279_g N_VSS_Mn9@2279_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2278 N_OUT9_Mn9@2278_d N_OUT8_Mn9@2278_g N_VSS_Mn9@2278_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2279 N_OUT9_Mp9@2279_d N_OUT8_Mp9@2279_g N_VDD_Mp9@2279_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2278 N_OUT9_Mp9@2278_d N_OUT8_Mp9@2278_g N_VDD_Mp9@2278_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2277 N_OUT9_Mn9@2277_d N_OUT8_Mn9@2277_g N_VSS_Mn9@2277_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2276 N_OUT9_Mn9@2276_d N_OUT8_Mn9@2276_g N_VSS_Mn9@2276_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2277 N_OUT9_Mp9@2277_d N_OUT8_Mp9@2277_g N_VDD_Mp9@2277_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2276 N_OUT9_Mp9@2276_d N_OUT8_Mp9@2276_g N_VDD_Mp9@2276_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2275 N_OUT9_Mn9@2275_d N_OUT8_Mn9@2275_g N_VSS_Mn9@2275_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2274 N_OUT9_Mn9@2274_d N_OUT8_Mn9@2274_g N_VSS_Mn9@2274_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2275 N_OUT9_Mp9@2275_d N_OUT8_Mp9@2275_g N_VDD_Mp9@2275_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2274 N_OUT9_Mp9@2274_d N_OUT8_Mp9@2274_g N_VDD_Mp9@2274_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2273 N_OUT9_Mn9@2273_d N_OUT8_Mn9@2273_g N_VSS_Mn9@2273_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2272 N_OUT9_Mn9@2272_d N_OUT8_Mn9@2272_g N_VSS_Mn9@2272_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2273 N_OUT9_Mp9@2273_d N_OUT8_Mp9@2273_g N_VDD_Mp9@2273_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2272 N_OUT9_Mp9@2272_d N_OUT8_Mp9@2272_g N_VDD_Mp9@2272_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2271 N_OUT9_Mn9@2271_d N_OUT8_Mn9@2271_g N_VSS_Mn9@2271_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2270 N_OUT9_Mn9@2270_d N_OUT8_Mn9@2270_g N_VSS_Mn9@2270_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2271 N_OUT9_Mp9@2271_d N_OUT8_Mp9@2271_g N_VDD_Mp9@2271_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2270 N_OUT9_Mp9@2270_d N_OUT8_Mp9@2270_g N_VDD_Mp9@2270_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2269 N_OUT9_Mn9@2269_d N_OUT8_Mn9@2269_g N_VSS_Mn9@2269_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2268 N_OUT9_Mn9@2268_d N_OUT8_Mn9@2268_g N_VSS_Mn9@2268_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2269 N_OUT9_Mp9@2269_d N_OUT8_Mp9@2269_g N_VDD_Mp9@2269_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2268 N_OUT9_Mp9@2268_d N_OUT8_Mp9@2268_g N_VDD_Mp9@2268_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2267 N_OUT9_Mn9@2267_d N_OUT8_Mn9@2267_g N_VSS_Mn9@2267_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2266 N_OUT9_Mn9@2266_d N_OUT8_Mn9@2266_g N_VSS_Mn9@2266_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2267 N_OUT9_Mp9@2267_d N_OUT8_Mp9@2267_g N_VDD_Mp9@2267_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2266 N_OUT9_Mp9@2266_d N_OUT8_Mp9@2266_g N_VDD_Mp9@2266_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2265 N_OUT9_Mn9@2265_d N_OUT8_Mn9@2265_g N_VSS_Mn9@2265_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2264 N_OUT9_Mn9@2264_d N_OUT8_Mn9@2264_g N_VSS_Mn9@2264_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2265 N_OUT9_Mp9@2265_d N_OUT8_Mp9@2265_g N_VDD_Mp9@2265_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2264 N_OUT9_Mp9@2264_d N_OUT8_Mp9@2264_g N_VDD_Mp9@2264_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2263 N_OUT9_Mn9@2263_d N_OUT8_Mn9@2263_g N_VSS_Mn9@2263_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2262 N_OUT9_Mn9@2262_d N_OUT8_Mn9@2262_g N_VSS_Mn9@2262_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2263 N_OUT9_Mp9@2263_d N_OUT8_Mp9@2263_g N_VDD_Mp9@2263_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2262 N_OUT9_Mp9@2262_d N_OUT8_Mp9@2262_g N_VDD_Mp9@2262_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2261 N_OUT9_Mn9@2261_d N_OUT8_Mn9@2261_g N_VSS_Mn9@2261_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2260 N_OUT9_Mn9@2260_d N_OUT8_Mn9@2260_g N_VSS_Mn9@2260_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2261 N_OUT9_Mp9@2261_d N_OUT8_Mp9@2261_g N_VDD_Mp9@2261_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2260 N_OUT9_Mp9@2260_d N_OUT8_Mp9@2260_g N_VDD_Mp9@2260_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2259 N_OUT9_Mn9@2259_d N_OUT8_Mn9@2259_g N_VSS_Mn9@2259_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2258 N_OUT9_Mn9@2258_d N_OUT8_Mn9@2258_g N_VSS_Mn9@2258_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2259 N_OUT9_Mp9@2259_d N_OUT8_Mp9@2259_g N_VDD_Mp9@2259_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2258 N_OUT9_Mp9@2258_d N_OUT8_Mp9@2258_g N_VDD_Mp9@2258_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2257 N_OUT9_Mn9@2257_d N_OUT8_Mn9@2257_g N_VSS_Mn9@2257_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2256 N_OUT9_Mn9@2256_d N_OUT8_Mn9@2256_g N_VSS_Mn9@2256_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2257 N_OUT9_Mp9@2257_d N_OUT8_Mp9@2257_g N_VDD_Mp9@2257_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2256 N_OUT9_Mp9@2256_d N_OUT8_Mp9@2256_g N_VDD_Mp9@2256_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2255 N_OUT9_Mn9@2255_d N_OUT8_Mn9@2255_g N_VSS_Mn9@2255_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2254 N_OUT9_Mn9@2254_d N_OUT8_Mn9@2254_g N_VSS_Mn9@2254_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2255 N_OUT9_Mp9@2255_d N_OUT8_Mp9@2255_g N_VDD_Mp9@2255_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2254 N_OUT9_Mp9@2254_d N_OUT8_Mp9@2254_g N_VDD_Mp9@2254_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2253 N_OUT9_Mn9@2253_d N_OUT8_Mn9@2253_g N_VSS_Mn9@2253_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2252 N_OUT9_Mn9@2252_d N_OUT8_Mn9@2252_g N_VSS_Mn9@2252_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2253 N_OUT9_Mp9@2253_d N_OUT8_Mp9@2253_g N_VDD_Mp9@2253_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2252 N_OUT9_Mp9@2252_d N_OUT8_Mp9@2252_g N_VDD_Mp9@2252_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2251 N_OUT9_Mn9@2251_d N_OUT8_Mn9@2251_g N_VSS_Mn9@2251_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2250 N_OUT9_Mn9@2250_d N_OUT8_Mn9@2250_g N_VSS_Mn9@2250_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2251 N_OUT9_Mp9@2251_d N_OUT8_Mp9@2251_g N_VDD_Mp9@2251_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2250 N_OUT9_Mp9@2250_d N_OUT8_Mp9@2250_g N_VDD_Mp9@2250_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2249 N_OUT9_Mn9@2249_d N_OUT8_Mn9@2249_g N_VSS_Mn9@2249_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2248 N_OUT9_Mn9@2248_d N_OUT8_Mn9@2248_g N_VSS_Mn9@2248_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2249 N_OUT9_Mp9@2249_d N_OUT8_Mp9@2249_g N_VDD_Mp9@2249_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2248 N_OUT9_Mp9@2248_d N_OUT8_Mp9@2248_g N_VDD_Mp9@2248_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2247 N_OUT9_Mn9@2247_d N_OUT8_Mn9@2247_g N_VSS_Mn9@2247_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2246 N_OUT9_Mn9@2246_d N_OUT8_Mn9@2246_g N_VSS_Mn9@2246_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2247 N_OUT9_Mp9@2247_d N_OUT8_Mp9@2247_g N_VDD_Mp9@2247_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2246 N_OUT9_Mp9@2246_d N_OUT8_Mp9@2246_g N_VDD_Mp9@2246_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2245 N_OUT9_Mn9@2245_d N_OUT8_Mn9@2245_g N_VSS_Mn9@2245_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2244 N_OUT9_Mn9@2244_d N_OUT8_Mn9@2244_g N_VSS_Mn9@2244_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2245 N_OUT9_Mp9@2245_d N_OUT8_Mp9@2245_g N_VDD_Mp9@2245_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2244 N_OUT9_Mp9@2244_d N_OUT8_Mp9@2244_g N_VDD_Mp9@2244_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2243 N_OUT9_Mn9@2243_d N_OUT8_Mn9@2243_g N_VSS_Mn9@2243_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2242 N_OUT9_Mn9@2242_d N_OUT8_Mn9@2242_g N_VSS_Mn9@2242_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2243 N_OUT9_Mp9@2243_d N_OUT8_Mp9@2243_g N_VDD_Mp9@2243_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2242 N_OUT9_Mp9@2242_d N_OUT8_Mp9@2242_g N_VDD_Mp9@2242_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2241 N_OUT9_Mn9@2241_d N_OUT8_Mn9@2241_g N_VSS_Mn9@2241_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2240 N_OUT9_Mn9@2240_d N_OUT8_Mn9@2240_g N_VSS_Mn9@2240_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2241 N_OUT9_Mp9@2241_d N_OUT8_Mp9@2241_g N_VDD_Mp9@2241_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2240 N_OUT9_Mp9@2240_d N_OUT8_Mp9@2240_g N_VDD_Mp9@2240_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2239 N_OUT9_Mn9@2239_d N_OUT8_Mn9@2239_g N_VSS_Mn9@2239_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2238 N_OUT9_Mn9@2238_d N_OUT8_Mn9@2238_g N_VSS_Mn9@2238_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2239 N_OUT9_Mp9@2239_d N_OUT8_Mp9@2239_g N_VDD_Mp9@2239_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2238 N_OUT9_Mp9@2238_d N_OUT8_Mp9@2238_g N_VDD_Mp9@2238_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2237 N_OUT9_Mn9@2237_d N_OUT8_Mn9@2237_g N_VSS_Mn9@2237_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2236 N_OUT9_Mn9@2236_d N_OUT8_Mn9@2236_g N_VSS_Mn9@2236_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2237 N_OUT9_Mp9@2237_d N_OUT8_Mp9@2237_g N_VDD_Mp9@2237_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2236 N_OUT9_Mp9@2236_d N_OUT8_Mp9@2236_g N_VDD_Mp9@2236_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2235 N_OUT9_Mn9@2235_d N_OUT8_Mn9@2235_g N_VSS_Mn9@2235_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2234 N_OUT9_Mn9@2234_d N_OUT8_Mn9@2234_g N_VSS_Mn9@2234_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2235 N_OUT9_Mp9@2235_d N_OUT8_Mp9@2235_g N_VDD_Mp9@2235_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2234 N_OUT9_Mp9@2234_d N_OUT8_Mp9@2234_g N_VDD_Mp9@2234_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2233 N_OUT9_Mn9@2233_d N_OUT8_Mn9@2233_g N_VSS_Mn9@2233_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2232 N_OUT9_Mn9@2232_d N_OUT8_Mn9@2232_g N_VSS_Mn9@2232_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2233 N_OUT9_Mp9@2233_d N_OUT8_Mp9@2233_g N_VDD_Mp9@2233_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2232 N_OUT9_Mp9@2232_d N_OUT8_Mp9@2232_g N_VDD_Mp9@2232_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2231 N_OUT9_Mn9@2231_d N_OUT8_Mn9@2231_g N_VSS_Mn9@2231_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2230 N_OUT9_Mn9@2230_d N_OUT8_Mn9@2230_g N_VSS_Mn9@2230_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2231 N_OUT9_Mp9@2231_d N_OUT8_Mp9@2231_g N_VDD_Mp9@2231_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2230 N_OUT9_Mp9@2230_d N_OUT8_Mp9@2230_g N_VDD_Mp9@2230_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2229 N_OUT9_Mn9@2229_d N_OUT8_Mn9@2229_g N_VSS_Mn9@2229_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2228 N_OUT9_Mn9@2228_d N_OUT8_Mn9@2228_g N_VSS_Mn9@2228_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2229 N_OUT9_Mp9@2229_d N_OUT8_Mp9@2229_g N_VDD_Mp9@2229_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2228 N_OUT9_Mp9@2228_d N_OUT8_Mp9@2228_g N_VDD_Mp9@2228_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2227 N_OUT9_Mn9@2227_d N_OUT8_Mn9@2227_g N_VSS_Mn9@2227_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2226 N_OUT9_Mn9@2226_d N_OUT8_Mn9@2226_g N_VSS_Mn9@2226_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2227 N_OUT9_Mp9@2227_d N_OUT8_Mp9@2227_g N_VDD_Mp9@2227_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2226 N_OUT9_Mp9@2226_d N_OUT8_Mp9@2226_g N_VDD_Mp9@2226_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2225 N_OUT9_Mn9@2225_d N_OUT8_Mn9@2225_g N_VSS_Mn9@2225_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2224 N_OUT9_Mn9@2224_d N_OUT8_Mn9@2224_g N_VSS_Mn9@2224_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2225 N_OUT9_Mp9@2225_d N_OUT8_Mp9@2225_g N_VDD_Mp9@2225_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2224 N_OUT9_Mp9@2224_d N_OUT8_Mp9@2224_g N_VDD_Mp9@2224_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2223 N_OUT9_Mn9@2223_d N_OUT8_Mn9@2223_g N_VSS_Mn9@2223_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2222 N_OUT9_Mn9@2222_d N_OUT8_Mn9@2222_g N_VSS_Mn9@2222_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2223 N_OUT9_Mp9@2223_d N_OUT8_Mp9@2223_g N_VDD_Mp9@2223_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2222 N_OUT9_Mp9@2222_d N_OUT8_Mp9@2222_g N_VDD_Mp9@2222_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2221 N_OUT9_Mn9@2221_d N_OUT8_Mn9@2221_g N_VSS_Mn9@2221_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2220 N_OUT9_Mn9@2220_d N_OUT8_Mn9@2220_g N_VSS_Mn9@2220_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2221 N_OUT9_Mp9@2221_d N_OUT8_Mp9@2221_g N_VDD_Mp9@2221_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2220 N_OUT9_Mp9@2220_d N_OUT8_Mp9@2220_g N_VDD_Mp9@2220_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2219 N_OUT9_Mn9@2219_d N_OUT8_Mn9@2219_g N_VSS_Mn9@2219_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2218 N_OUT9_Mn9@2218_d N_OUT8_Mn9@2218_g N_VSS_Mn9@2218_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2219 N_OUT9_Mp9@2219_d N_OUT8_Mp9@2219_g N_VDD_Mp9@2219_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2218 N_OUT9_Mp9@2218_d N_OUT8_Mp9@2218_g N_VDD_Mp9@2218_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2217 N_OUT9_Mn9@2217_d N_OUT8_Mn9@2217_g N_VSS_Mn9@2217_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2216 N_OUT9_Mn9@2216_d N_OUT8_Mn9@2216_g N_VSS_Mn9@2216_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2217 N_OUT9_Mp9@2217_d N_OUT8_Mp9@2217_g N_VDD_Mp9@2217_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2216 N_OUT9_Mp9@2216_d N_OUT8_Mp9@2216_g N_VDD_Mp9@2216_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2215 N_OUT9_Mn9@2215_d N_OUT8_Mn9@2215_g N_VSS_Mn9@2215_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2214 N_OUT9_Mn9@2214_d N_OUT8_Mn9@2214_g N_VSS_Mn9@2214_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2215 N_OUT9_Mp9@2215_d N_OUT8_Mp9@2215_g N_VDD_Mp9@2215_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2214 N_OUT9_Mp9@2214_d N_OUT8_Mp9@2214_g N_VDD_Mp9@2214_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2213 N_OUT9_Mn9@2213_d N_OUT8_Mn9@2213_g N_VSS_Mn9@2213_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2212 N_OUT9_Mn9@2212_d N_OUT8_Mn9@2212_g N_VSS_Mn9@2212_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2213 N_OUT9_Mp9@2213_d N_OUT8_Mp9@2213_g N_VDD_Mp9@2213_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2212 N_OUT9_Mp9@2212_d N_OUT8_Mp9@2212_g N_VDD_Mp9@2212_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2211 N_OUT9_Mn9@2211_d N_OUT8_Mn9@2211_g N_VSS_Mn9@2211_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2210 N_OUT9_Mn9@2210_d N_OUT8_Mn9@2210_g N_VSS_Mn9@2210_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2211 N_OUT9_Mp9@2211_d N_OUT8_Mp9@2211_g N_VDD_Mp9@2211_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2210 N_OUT9_Mp9@2210_d N_OUT8_Mp9@2210_g N_VDD_Mp9@2210_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2209 N_OUT9_Mn9@2209_d N_OUT8_Mn9@2209_g N_VSS_Mn9@2209_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2208 N_OUT9_Mn9@2208_d N_OUT8_Mn9@2208_g N_VSS_Mn9@2208_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2209 N_OUT9_Mp9@2209_d N_OUT8_Mp9@2209_g N_VDD_Mp9@2209_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2208 N_OUT9_Mp9@2208_d N_OUT8_Mp9@2208_g N_VDD_Mp9@2208_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2207 N_OUT9_Mn9@2207_d N_OUT8_Mn9@2207_g N_VSS_Mn9@2207_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2206 N_OUT9_Mn9@2206_d N_OUT8_Mn9@2206_g N_VSS_Mn9@2206_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2207 N_OUT9_Mp9@2207_d N_OUT8_Mp9@2207_g N_VDD_Mp9@2207_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2206 N_OUT9_Mp9@2206_d N_OUT8_Mp9@2206_g N_VDD_Mp9@2206_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2205 N_OUT9_Mn9@2205_d N_OUT8_Mn9@2205_g N_VSS_Mn9@2205_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2204 N_OUT9_Mn9@2204_d N_OUT8_Mn9@2204_g N_VSS_Mn9@2204_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2205 N_OUT9_Mp9@2205_d N_OUT8_Mp9@2205_g N_VDD_Mp9@2205_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2204 N_OUT9_Mp9@2204_d N_OUT8_Mp9@2204_g N_VDD_Mp9@2204_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2203 N_OUT9_Mn9@2203_d N_OUT8_Mn9@2203_g N_VSS_Mn9@2203_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2202 N_OUT9_Mn9@2202_d N_OUT8_Mn9@2202_g N_VSS_Mn9@2202_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2203 N_OUT9_Mp9@2203_d N_OUT8_Mp9@2203_g N_VDD_Mp9@2203_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2202 N_OUT9_Mp9@2202_d N_OUT8_Mp9@2202_g N_VDD_Mp9@2202_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2201 N_OUT9_Mn9@2201_d N_OUT8_Mn9@2201_g N_VSS_Mn9@2201_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2200 N_OUT9_Mn9@2200_d N_OUT8_Mn9@2200_g N_VSS_Mn9@2200_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2201 N_OUT9_Mp9@2201_d N_OUT8_Mp9@2201_g N_VDD_Mp9@2201_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2200 N_OUT9_Mp9@2200_d N_OUT8_Mp9@2200_g N_VDD_Mp9@2200_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2199 N_OUT9_Mn9@2199_d N_OUT8_Mn9@2199_g N_VSS_Mn9@2199_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2198 N_OUT9_Mn9@2198_d N_OUT8_Mn9@2198_g N_VSS_Mn9@2198_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2199 N_OUT9_Mp9@2199_d N_OUT8_Mp9@2199_g N_VDD_Mp9@2199_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2198 N_OUT9_Mp9@2198_d N_OUT8_Mp9@2198_g N_VDD_Mp9@2198_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2197 N_OUT9_Mn9@2197_d N_OUT8_Mn9@2197_g N_VSS_Mn9@2197_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2196 N_OUT9_Mn9@2196_d N_OUT8_Mn9@2196_g N_VSS_Mn9@2196_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2197 N_OUT9_Mp9@2197_d N_OUT8_Mp9@2197_g N_VDD_Mp9@2197_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2196 N_OUT9_Mp9@2196_d N_OUT8_Mp9@2196_g N_VDD_Mp9@2196_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2195 N_OUT9_Mn9@2195_d N_OUT8_Mn9@2195_g N_VSS_Mn9@2195_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2194 N_OUT9_Mn9@2194_d N_OUT8_Mn9@2194_g N_VSS_Mn9@2194_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2195 N_OUT9_Mp9@2195_d N_OUT8_Mp9@2195_g N_VDD_Mp9@2195_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2194 N_OUT9_Mp9@2194_d N_OUT8_Mp9@2194_g N_VDD_Mp9@2194_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2193 N_OUT9_Mn9@2193_d N_OUT8_Mn9@2193_g N_VSS_Mn9@2193_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2192 N_OUT9_Mn9@2192_d N_OUT8_Mn9@2192_g N_VSS_Mn9@2192_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2193 N_OUT9_Mp9@2193_d N_OUT8_Mp9@2193_g N_VDD_Mp9@2193_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2192 N_OUT9_Mp9@2192_d N_OUT8_Mp9@2192_g N_VDD_Mp9@2192_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2191 N_OUT9_Mn9@2191_d N_OUT8_Mn9@2191_g N_VSS_Mn9@2191_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2190 N_OUT9_Mn9@2190_d N_OUT8_Mn9@2190_g N_VSS_Mn9@2190_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2191 N_OUT9_Mp9@2191_d N_OUT8_Mp9@2191_g N_VDD_Mp9@2191_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2190 N_OUT9_Mp9@2190_d N_OUT8_Mp9@2190_g N_VDD_Mp9@2190_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2189 N_OUT9_Mn9@2189_d N_OUT8_Mn9@2189_g N_VSS_Mn9@2189_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2188 N_OUT9_Mn9@2188_d N_OUT8_Mn9@2188_g N_VSS_Mn9@2188_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2189 N_OUT9_Mp9@2189_d N_OUT8_Mp9@2189_g N_VDD_Mp9@2189_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2188 N_OUT9_Mp9@2188_d N_OUT8_Mp9@2188_g N_VDD_Mp9@2188_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2187 N_OUT9_Mn9@2187_d N_OUT8_Mn9@2187_g N_VSS_Mn9@2187_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2186 N_OUT9_Mn9@2186_d N_OUT8_Mn9@2186_g N_VSS_Mn9@2186_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2187 N_OUT9_Mp9@2187_d N_OUT8_Mp9@2187_g N_VDD_Mp9@2187_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2186 N_OUT9_Mp9@2186_d N_OUT8_Mp9@2186_g N_VDD_Mp9@2186_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2185 N_OUT9_Mn9@2185_d N_OUT8_Mn9@2185_g N_VSS_Mn9@2185_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2184 N_OUT9_Mn9@2184_d N_OUT8_Mn9@2184_g N_VSS_Mn9@2184_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2185 N_OUT9_Mp9@2185_d N_OUT8_Mp9@2185_g N_VDD_Mp9@2185_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2184 N_OUT9_Mp9@2184_d N_OUT8_Mp9@2184_g N_VDD_Mp9@2184_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2183 N_OUT9_Mn9@2183_d N_OUT8_Mn9@2183_g N_VSS_Mn9@2183_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2182 N_OUT9_Mn9@2182_d N_OUT8_Mn9@2182_g N_VSS_Mn9@2182_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2183 N_OUT9_Mp9@2183_d N_OUT8_Mp9@2183_g N_VDD_Mp9@2183_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2182 N_OUT9_Mp9@2182_d N_OUT8_Mp9@2182_g N_VDD_Mp9@2182_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2181 N_OUT9_Mn9@2181_d N_OUT8_Mn9@2181_g N_VSS_Mn9@2181_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2180 N_OUT9_Mn9@2180_d N_OUT8_Mn9@2180_g N_VSS_Mn9@2180_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2181 N_OUT9_Mp9@2181_d N_OUT8_Mp9@2181_g N_VDD_Mp9@2181_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2180 N_OUT9_Mp9@2180_d N_OUT8_Mp9@2180_g N_VDD_Mp9@2180_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2179 N_OUT9_Mn9@2179_d N_OUT8_Mn9@2179_g N_VSS_Mn9@2179_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2178 N_OUT9_Mn9@2178_d N_OUT8_Mn9@2178_g N_VSS_Mn9@2178_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2179 N_OUT9_Mp9@2179_d N_OUT8_Mp9@2179_g N_VDD_Mp9@2179_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2178 N_OUT9_Mp9@2178_d N_OUT8_Mp9@2178_g N_VDD_Mp9@2178_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2177 N_OUT9_Mn9@2177_d N_OUT8_Mn9@2177_g N_VSS_Mn9@2177_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2176 N_OUT9_Mn9@2176_d N_OUT8_Mn9@2176_g N_VSS_Mn9@2176_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2177 N_OUT9_Mp9@2177_d N_OUT8_Mp9@2177_g N_VDD_Mp9@2177_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2176 N_OUT9_Mp9@2176_d N_OUT8_Mp9@2176_g N_VDD_Mp9@2176_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2175 N_OUT9_Mn9@2175_d N_OUT8_Mn9@2175_g N_VSS_Mn9@2175_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2174 N_OUT9_Mn9@2174_d N_OUT8_Mn9@2174_g N_VSS_Mn9@2174_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2175 N_OUT9_Mp9@2175_d N_OUT8_Mp9@2175_g N_VDD_Mp9@2175_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2174 N_OUT9_Mp9@2174_d N_OUT8_Mp9@2174_g N_VDD_Mp9@2174_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2173 N_OUT9_Mn9@2173_d N_OUT8_Mn9@2173_g N_VSS_Mn9@2173_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2172 N_OUT9_Mn9@2172_d N_OUT8_Mn9@2172_g N_VSS_Mn9@2172_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2173 N_OUT9_Mp9@2173_d N_OUT8_Mp9@2173_g N_VDD_Mp9@2173_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2172 N_OUT9_Mp9@2172_d N_OUT8_Mp9@2172_g N_VDD_Mp9@2172_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2171 N_OUT9_Mn9@2171_d N_OUT8_Mn9@2171_g N_VSS_Mn9@2171_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2170 N_OUT9_Mn9@2170_d N_OUT8_Mn9@2170_g N_VSS_Mn9@2170_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2171 N_OUT9_Mp9@2171_d N_OUT8_Mp9@2171_g N_VDD_Mp9@2171_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2170 N_OUT9_Mp9@2170_d N_OUT8_Mp9@2170_g N_VDD_Mp9@2170_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2169 N_OUT9_Mn9@2169_d N_OUT8_Mn9@2169_g N_VSS_Mn9@2169_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2168 N_OUT9_Mn9@2168_d N_OUT8_Mn9@2168_g N_VSS_Mn9@2168_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2169 N_OUT9_Mp9@2169_d N_OUT8_Mp9@2169_g N_VDD_Mp9@2169_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2168 N_OUT9_Mp9@2168_d N_OUT8_Mp9@2168_g N_VDD_Mp9@2168_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2167 N_OUT9_Mn9@2167_d N_OUT8_Mn9@2167_g N_VSS_Mn9@2167_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2166 N_OUT9_Mn9@2166_d N_OUT8_Mn9@2166_g N_VSS_Mn9@2166_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2167 N_OUT9_Mp9@2167_d N_OUT8_Mp9@2167_g N_VDD_Mp9@2167_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2166 N_OUT9_Mp9@2166_d N_OUT8_Mp9@2166_g N_VDD_Mp9@2166_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2165 N_OUT9_Mn9@2165_d N_OUT8_Mn9@2165_g N_VSS_Mn9@2165_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2164 N_OUT9_Mn9@2164_d N_OUT8_Mn9@2164_g N_VSS_Mn9@2164_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2165 N_OUT9_Mp9@2165_d N_OUT8_Mp9@2165_g N_VDD_Mp9@2165_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2164 N_OUT9_Mp9@2164_d N_OUT8_Mp9@2164_g N_VDD_Mp9@2164_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2163 N_OUT9_Mn9@2163_d N_OUT8_Mn9@2163_g N_VSS_Mn9@2163_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2162 N_OUT9_Mn9@2162_d N_OUT8_Mn9@2162_g N_VSS_Mn9@2162_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2163 N_OUT9_Mp9@2163_d N_OUT8_Mp9@2163_g N_VDD_Mp9@2163_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2162 N_OUT9_Mp9@2162_d N_OUT8_Mp9@2162_g N_VDD_Mp9@2162_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2161 N_OUT9_Mn9@2161_d N_OUT8_Mn9@2161_g N_VSS_Mn9@2161_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2160 N_OUT9_Mn9@2160_d N_OUT8_Mn9@2160_g N_VSS_Mn9@2160_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2161 N_OUT9_Mp9@2161_d N_OUT8_Mp9@2161_g N_VDD_Mp9@2161_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2160 N_OUT9_Mp9@2160_d N_OUT8_Mp9@2160_g N_VDD_Mp9@2160_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2159 N_OUT9_Mn9@2159_d N_OUT8_Mn9@2159_g N_VSS_Mn9@2159_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2158 N_OUT9_Mn9@2158_d N_OUT8_Mn9@2158_g N_VSS_Mn9@2158_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2159 N_OUT9_Mp9@2159_d N_OUT8_Mp9@2159_g N_VDD_Mp9@2159_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2158 N_OUT9_Mp9@2158_d N_OUT8_Mp9@2158_g N_VDD_Mp9@2158_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2157 N_OUT9_Mn9@2157_d N_OUT8_Mn9@2157_g N_VSS_Mn9@2157_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2156 N_OUT9_Mn9@2156_d N_OUT8_Mn9@2156_g N_VSS_Mn9@2156_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2157 N_OUT9_Mp9@2157_d N_OUT8_Mp9@2157_g N_VDD_Mp9@2157_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2156 N_OUT9_Mp9@2156_d N_OUT8_Mp9@2156_g N_VDD_Mp9@2156_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2155 N_OUT9_Mn9@2155_d N_OUT8_Mn9@2155_g N_VSS_Mn9@2155_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2154 N_OUT9_Mn9@2154_d N_OUT8_Mn9@2154_g N_VSS_Mn9@2154_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2155 N_OUT9_Mp9@2155_d N_OUT8_Mp9@2155_g N_VDD_Mp9@2155_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2154 N_OUT9_Mp9@2154_d N_OUT8_Mp9@2154_g N_VDD_Mp9@2154_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2153 N_OUT9_Mn9@2153_d N_OUT8_Mn9@2153_g N_VSS_Mn9@2153_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2152 N_OUT9_Mn9@2152_d N_OUT8_Mn9@2152_g N_VSS_Mn9@2152_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2153 N_OUT9_Mp9@2153_d N_OUT8_Mp9@2153_g N_VDD_Mp9@2153_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2152 N_OUT9_Mp9@2152_d N_OUT8_Mp9@2152_g N_VDD_Mp9@2152_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2151 N_OUT9_Mn9@2151_d N_OUT8_Mn9@2151_g N_VSS_Mn9@2151_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2150 N_OUT9_Mn9@2150_d N_OUT8_Mn9@2150_g N_VSS_Mn9@2150_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2151 N_OUT9_Mp9@2151_d N_OUT8_Mp9@2151_g N_VDD_Mp9@2151_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2150 N_OUT9_Mp9@2150_d N_OUT8_Mp9@2150_g N_VDD_Mp9@2150_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2149 N_OUT9_Mn9@2149_d N_OUT8_Mn9@2149_g N_VSS_Mn9@2149_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2148 N_OUT9_Mn9@2148_d N_OUT8_Mn9@2148_g N_VSS_Mn9@2148_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2149 N_OUT9_Mp9@2149_d N_OUT8_Mp9@2149_g N_VDD_Mp9@2149_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2148 N_OUT9_Mp9@2148_d N_OUT8_Mp9@2148_g N_VDD_Mp9@2148_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2147 N_OUT9_Mn9@2147_d N_OUT8_Mn9@2147_g N_VSS_Mn9@2147_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2146 N_OUT9_Mn9@2146_d N_OUT8_Mn9@2146_g N_VSS_Mn9@2146_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2147 N_OUT9_Mp9@2147_d N_OUT8_Mp9@2147_g N_VDD_Mp9@2147_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2146 N_OUT9_Mp9@2146_d N_OUT8_Mp9@2146_g N_VDD_Mp9@2146_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2145 N_OUT9_Mn9@2145_d N_OUT8_Mn9@2145_g N_VSS_Mn9@2145_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2144 N_OUT9_Mn9@2144_d N_OUT8_Mn9@2144_g N_VSS_Mn9@2144_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2145 N_OUT9_Mp9@2145_d N_OUT8_Mp9@2145_g N_VDD_Mp9@2145_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2144 N_OUT9_Mp9@2144_d N_OUT8_Mp9@2144_g N_VDD_Mp9@2144_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2143 N_OUT9_Mn9@2143_d N_OUT8_Mn9@2143_g N_VSS_Mn9@2143_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2142 N_OUT9_Mn9@2142_d N_OUT8_Mn9@2142_g N_VSS_Mn9@2142_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2143 N_OUT9_Mp9@2143_d N_OUT8_Mp9@2143_g N_VDD_Mp9@2143_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2142 N_OUT9_Mp9@2142_d N_OUT8_Mp9@2142_g N_VDD_Mp9@2142_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2141 N_OUT9_Mn9@2141_d N_OUT8_Mn9@2141_g N_VSS_Mn9@2141_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2140 N_OUT9_Mn9@2140_d N_OUT8_Mn9@2140_g N_VSS_Mn9@2140_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2141 N_OUT9_Mp9@2141_d N_OUT8_Mp9@2141_g N_VDD_Mp9@2141_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2140 N_OUT9_Mp9@2140_d N_OUT8_Mp9@2140_g N_VDD_Mp9@2140_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2139 N_OUT9_Mn9@2139_d N_OUT8_Mn9@2139_g N_VSS_Mn9@2139_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2138 N_OUT9_Mn9@2138_d N_OUT8_Mn9@2138_g N_VSS_Mn9@2138_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2139 N_OUT9_Mp9@2139_d N_OUT8_Mp9@2139_g N_VDD_Mp9@2139_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2138 N_OUT9_Mp9@2138_d N_OUT8_Mp9@2138_g N_VDD_Mp9@2138_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2137 N_OUT9_Mn9@2137_d N_OUT8_Mn9@2137_g N_VSS_Mn9@2137_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2136 N_OUT9_Mn9@2136_d N_OUT8_Mn9@2136_g N_VSS_Mn9@2136_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2137 N_OUT9_Mp9@2137_d N_OUT8_Mp9@2137_g N_VDD_Mp9@2137_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2136 N_OUT9_Mp9@2136_d N_OUT8_Mp9@2136_g N_VDD_Mp9@2136_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2135 N_OUT9_Mn9@2135_d N_OUT8_Mn9@2135_g N_VSS_Mn9@2135_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2134 N_OUT9_Mn9@2134_d N_OUT8_Mn9@2134_g N_VSS_Mn9@2134_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2135 N_OUT9_Mp9@2135_d N_OUT8_Mp9@2135_g N_VDD_Mp9@2135_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2134 N_OUT9_Mp9@2134_d N_OUT8_Mp9@2134_g N_VDD_Mp9@2134_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2133 N_OUT9_Mn9@2133_d N_OUT8_Mn9@2133_g N_VSS_Mn9@2133_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2132 N_OUT9_Mn9@2132_d N_OUT8_Mn9@2132_g N_VSS_Mn9@2132_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2133 N_OUT9_Mp9@2133_d N_OUT8_Mp9@2133_g N_VDD_Mp9@2133_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2132 N_OUT9_Mp9@2132_d N_OUT8_Mp9@2132_g N_VDD_Mp9@2132_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2131 N_OUT9_Mn9@2131_d N_OUT8_Mn9@2131_g N_VSS_Mn9@2131_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2130 N_OUT9_Mn9@2130_d N_OUT8_Mn9@2130_g N_VSS_Mn9@2130_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2131 N_OUT9_Mp9@2131_d N_OUT8_Mp9@2131_g N_VDD_Mp9@2131_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2130 N_OUT9_Mp9@2130_d N_OUT8_Mp9@2130_g N_VDD_Mp9@2130_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2129 N_OUT9_Mn9@2129_d N_OUT8_Mn9@2129_g N_VSS_Mn9@2129_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2128 N_OUT9_Mn9@2128_d N_OUT8_Mn9@2128_g N_VSS_Mn9@2128_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2129 N_OUT9_Mp9@2129_d N_OUT8_Mp9@2129_g N_VDD_Mp9@2129_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2128 N_OUT9_Mp9@2128_d N_OUT8_Mp9@2128_g N_VDD_Mp9@2128_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2127 N_OUT9_Mn9@2127_d N_OUT8_Mn9@2127_g N_VSS_Mn9@2127_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2126 N_OUT9_Mn9@2126_d N_OUT8_Mn9@2126_g N_VSS_Mn9@2126_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2127 N_OUT9_Mp9@2127_d N_OUT8_Mp9@2127_g N_VDD_Mp9@2127_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2126 N_OUT9_Mp9@2126_d N_OUT8_Mp9@2126_g N_VDD_Mp9@2126_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2125 N_OUT9_Mn9@2125_d N_OUT8_Mn9@2125_g N_VSS_Mn9@2125_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2124 N_OUT9_Mn9@2124_d N_OUT8_Mn9@2124_g N_VSS_Mn9@2124_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2125 N_OUT9_Mp9@2125_d N_OUT8_Mp9@2125_g N_VDD_Mp9@2125_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2124 N_OUT9_Mp9@2124_d N_OUT8_Mp9@2124_g N_VDD_Mp9@2124_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2123 N_OUT9_Mn9@2123_d N_OUT8_Mn9@2123_g N_VSS_Mn9@2123_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2122 N_OUT9_Mn9@2122_d N_OUT8_Mn9@2122_g N_VSS_Mn9@2122_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2123 N_OUT9_Mp9@2123_d N_OUT8_Mp9@2123_g N_VDD_Mp9@2123_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2122 N_OUT9_Mp9@2122_d N_OUT8_Mp9@2122_g N_VDD_Mp9@2122_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2121 N_OUT9_Mn9@2121_d N_OUT8_Mn9@2121_g N_VSS_Mn9@2121_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2120 N_OUT9_Mn9@2120_d N_OUT8_Mn9@2120_g N_VSS_Mn9@2120_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2121 N_OUT9_Mp9@2121_d N_OUT8_Mp9@2121_g N_VDD_Mp9@2121_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2120 N_OUT9_Mp9@2120_d N_OUT8_Mp9@2120_g N_VDD_Mp9@2120_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2119 N_OUT9_Mn9@2119_d N_OUT8_Mn9@2119_g N_VSS_Mn9@2119_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2118 N_OUT9_Mn9@2118_d N_OUT8_Mn9@2118_g N_VSS_Mn9@2118_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2119 N_OUT9_Mp9@2119_d N_OUT8_Mp9@2119_g N_VDD_Mp9@2119_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2118 N_OUT9_Mp9@2118_d N_OUT8_Mp9@2118_g N_VDD_Mp9@2118_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2117 N_OUT9_Mn9@2117_d N_OUT8_Mn9@2117_g N_VSS_Mn9@2117_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2116 N_OUT9_Mn9@2116_d N_OUT8_Mn9@2116_g N_VSS_Mn9@2116_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2117 N_OUT9_Mp9@2117_d N_OUT8_Mp9@2117_g N_VDD_Mp9@2117_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2116 N_OUT9_Mp9@2116_d N_OUT8_Mp9@2116_g N_VDD_Mp9@2116_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2115 N_OUT9_Mn9@2115_d N_OUT8_Mn9@2115_g N_VSS_Mn9@2115_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2114 N_OUT9_Mn9@2114_d N_OUT8_Mn9@2114_g N_VSS_Mn9@2114_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2115 N_OUT9_Mp9@2115_d N_OUT8_Mp9@2115_g N_VDD_Mp9@2115_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2114 N_OUT9_Mp9@2114_d N_OUT8_Mp9@2114_g N_VDD_Mp9@2114_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2113 N_OUT9_Mn9@2113_d N_OUT8_Mn9@2113_g N_VSS_Mn9@2113_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2112 N_OUT9_Mn9@2112_d N_OUT8_Mn9@2112_g N_VSS_Mn9@2112_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2113 N_OUT9_Mp9@2113_d N_OUT8_Mp9@2113_g N_VDD_Mp9@2113_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2112 N_OUT9_Mp9@2112_d N_OUT8_Mp9@2112_g N_VDD_Mp9@2112_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2111 N_OUT9_Mn9@2111_d N_OUT8_Mn9@2111_g N_VSS_Mn9@2111_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2110 N_OUT9_Mn9@2110_d N_OUT8_Mn9@2110_g N_VSS_Mn9@2110_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2111 N_OUT9_Mp9@2111_d N_OUT8_Mp9@2111_g N_VDD_Mp9@2111_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2110 N_OUT9_Mp9@2110_d N_OUT8_Mp9@2110_g N_VDD_Mp9@2110_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2109 N_OUT9_Mn9@2109_d N_OUT8_Mn9@2109_g N_VSS_Mn9@2109_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2108 N_OUT9_Mn9@2108_d N_OUT8_Mn9@2108_g N_VSS_Mn9@2108_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2109 N_OUT9_Mp9@2109_d N_OUT8_Mp9@2109_g N_VDD_Mp9@2109_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2108 N_OUT9_Mp9@2108_d N_OUT8_Mp9@2108_g N_VDD_Mp9@2108_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2107 N_OUT9_Mn9@2107_d N_OUT8_Mn9@2107_g N_VSS_Mn9@2107_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2106 N_OUT9_Mn9@2106_d N_OUT8_Mn9@2106_g N_VSS_Mn9@2106_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2107 N_OUT9_Mp9@2107_d N_OUT8_Mp9@2107_g N_VDD_Mp9@2107_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2106 N_OUT9_Mp9@2106_d N_OUT8_Mp9@2106_g N_VDD_Mp9@2106_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2105 N_OUT9_Mn9@2105_d N_OUT8_Mn9@2105_g N_VSS_Mn9@2105_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2104 N_OUT9_Mn9@2104_d N_OUT8_Mn9@2104_g N_VSS_Mn9@2104_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2105 N_OUT9_Mp9@2105_d N_OUT8_Mp9@2105_g N_VDD_Mp9@2105_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2104 N_OUT9_Mp9@2104_d N_OUT8_Mp9@2104_g N_VDD_Mp9@2104_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2103 N_OUT9_Mn9@2103_d N_OUT8_Mn9@2103_g N_VSS_Mn9@2103_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2102 N_OUT9_Mn9@2102_d N_OUT8_Mn9@2102_g N_VSS_Mn9@2102_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2103 N_OUT9_Mp9@2103_d N_OUT8_Mp9@2103_g N_VDD_Mp9@2103_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2102 N_OUT9_Mp9@2102_d N_OUT8_Mp9@2102_g N_VDD_Mp9@2102_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2101 N_OUT9_Mn9@2101_d N_OUT8_Mn9@2101_g N_VSS_Mn9@2101_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2100 N_OUT9_Mn9@2100_d N_OUT8_Mn9@2100_g N_VSS_Mn9@2100_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2101 N_OUT9_Mp9@2101_d N_OUT8_Mp9@2101_g N_VDD_Mp9@2101_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2100 N_OUT9_Mp9@2100_d N_OUT8_Mp9@2100_g N_VDD_Mp9@2100_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2099 N_OUT9_Mn9@2099_d N_OUT8_Mn9@2099_g N_VSS_Mn9@2099_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2098 N_OUT9_Mn9@2098_d N_OUT8_Mn9@2098_g N_VSS_Mn9@2098_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2099 N_OUT9_Mp9@2099_d N_OUT8_Mp9@2099_g N_VDD_Mp9@2099_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2098 N_OUT9_Mp9@2098_d N_OUT8_Mp9@2098_g N_VDD_Mp9@2098_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2097 N_OUT9_Mn9@2097_d N_OUT8_Mn9@2097_g N_VSS_Mn9@2097_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2096 N_OUT9_Mn9@2096_d N_OUT8_Mn9@2096_g N_VSS_Mn9@2096_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2097 N_OUT9_Mp9@2097_d N_OUT8_Mp9@2097_g N_VDD_Mp9@2097_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2096 N_OUT9_Mp9@2096_d N_OUT8_Mp9@2096_g N_VDD_Mp9@2096_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2095 N_OUT9_Mn9@2095_d N_OUT8_Mn9@2095_g N_VSS_Mn9@2095_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2094 N_OUT9_Mn9@2094_d N_OUT8_Mn9@2094_g N_VSS_Mn9@2094_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2095 N_OUT9_Mp9@2095_d N_OUT8_Mp9@2095_g N_VDD_Mp9@2095_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2094 N_OUT9_Mp9@2094_d N_OUT8_Mp9@2094_g N_VDD_Mp9@2094_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2093 N_OUT9_Mn9@2093_d N_OUT8_Mn9@2093_g N_VSS_Mn9@2093_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2092 N_OUT9_Mn9@2092_d N_OUT8_Mn9@2092_g N_VSS_Mn9@2092_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2093 N_OUT9_Mp9@2093_d N_OUT8_Mp9@2093_g N_VDD_Mp9@2093_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2092 N_OUT9_Mp9@2092_d N_OUT8_Mp9@2092_g N_VDD_Mp9@2092_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2091 N_OUT9_Mn9@2091_d N_OUT8_Mn9@2091_g N_VSS_Mn9@2091_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2090 N_OUT9_Mn9@2090_d N_OUT8_Mn9@2090_g N_VSS_Mn9@2090_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2091 N_OUT9_Mp9@2091_d N_OUT8_Mp9@2091_g N_VDD_Mp9@2091_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2090 N_OUT9_Mp9@2090_d N_OUT8_Mp9@2090_g N_VDD_Mp9@2090_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2089 N_OUT9_Mn9@2089_d N_OUT8_Mn9@2089_g N_VSS_Mn9@2089_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2088 N_OUT9_Mn9@2088_d N_OUT8_Mn9@2088_g N_VSS_Mn9@2088_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2089 N_OUT9_Mp9@2089_d N_OUT8_Mp9@2089_g N_VDD_Mp9@2089_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2088 N_OUT9_Mp9@2088_d N_OUT8_Mp9@2088_g N_VDD_Mp9@2088_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2087 N_OUT9_Mn9@2087_d N_OUT8_Mn9@2087_g N_VSS_Mn9@2087_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2086 N_OUT9_Mn9@2086_d N_OUT8_Mn9@2086_g N_VSS_Mn9@2086_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2087 N_OUT9_Mp9@2087_d N_OUT8_Mp9@2087_g N_VDD_Mp9@2087_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2086 N_OUT9_Mp9@2086_d N_OUT8_Mp9@2086_g N_VDD_Mp9@2086_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2085 N_OUT9_Mn9@2085_d N_OUT8_Mn9@2085_g N_VSS_Mn9@2085_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2084 N_OUT9_Mn9@2084_d N_OUT8_Mn9@2084_g N_VSS_Mn9@2084_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2085 N_OUT9_Mp9@2085_d N_OUT8_Mp9@2085_g N_VDD_Mp9@2085_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2084 N_OUT9_Mp9@2084_d N_OUT8_Mp9@2084_g N_VDD_Mp9@2084_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2083 N_OUT9_Mn9@2083_d N_OUT8_Mn9@2083_g N_VSS_Mn9@2083_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2082 N_OUT9_Mn9@2082_d N_OUT8_Mn9@2082_g N_VSS_Mn9@2082_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2083 N_OUT9_Mp9@2083_d N_OUT8_Mp9@2083_g N_VDD_Mp9@2083_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2082 N_OUT9_Mp9@2082_d N_OUT8_Mp9@2082_g N_VDD_Mp9@2082_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2081 N_OUT9_Mn9@2081_d N_OUT8_Mn9@2081_g N_VSS_Mn9@2081_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2080 N_OUT9_Mn9@2080_d N_OUT8_Mn9@2080_g N_VSS_Mn9@2080_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2081 N_OUT9_Mp9@2081_d N_OUT8_Mp9@2081_g N_VDD_Mp9@2081_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2080 N_OUT9_Mp9@2080_d N_OUT8_Mp9@2080_g N_VDD_Mp9@2080_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2079 N_OUT9_Mn9@2079_d N_OUT8_Mn9@2079_g N_VSS_Mn9@2079_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2078 N_OUT9_Mn9@2078_d N_OUT8_Mn9@2078_g N_VSS_Mn9@2078_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2079 N_OUT9_Mp9@2079_d N_OUT8_Mp9@2079_g N_VDD_Mp9@2079_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2078 N_OUT9_Mp9@2078_d N_OUT8_Mp9@2078_g N_VDD_Mp9@2078_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2077 N_OUT9_Mn9@2077_d N_OUT8_Mn9@2077_g N_VSS_Mn9@2077_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2076 N_OUT9_Mn9@2076_d N_OUT8_Mn9@2076_g N_VSS_Mn9@2076_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2077 N_OUT9_Mp9@2077_d N_OUT8_Mp9@2077_g N_VDD_Mp9@2077_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2076 N_OUT9_Mp9@2076_d N_OUT8_Mp9@2076_g N_VDD_Mp9@2076_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2075 N_OUT9_Mn9@2075_d N_OUT8_Mn9@2075_g N_VSS_Mn9@2075_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2074 N_OUT9_Mn9@2074_d N_OUT8_Mn9@2074_g N_VSS_Mn9@2074_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2075 N_OUT9_Mp9@2075_d N_OUT8_Mp9@2075_g N_VDD_Mp9@2075_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2074 N_OUT9_Mp9@2074_d N_OUT8_Mp9@2074_g N_VDD_Mp9@2074_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2073 N_OUT9_Mn9@2073_d N_OUT8_Mn9@2073_g N_VSS_Mn9@2073_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2072 N_OUT9_Mn9@2072_d N_OUT8_Mn9@2072_g N_VSS_Mn9@2072_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2073 N_OUT9_Mp9@2073_d N_OUT8_Mp9@2073_g N_VDD_Mp9@2073_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2072 N_OUT9_Mp9@2072_d N_OUT8_Mp9@2072_g N_VDD_Mp9@2072_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2071 N_OUT9_Mn9@2071_d N_OUT8_Mn9@2071_g N_VSS_Mn9@2071_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2070 N_OUT9_Mn9@2070_d N_OUT8_Mn9@2070_g N_VSS_Mn9@2070_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2071 N_OUT9_Mp9@2071_d N_OUT8_Mp9@2071_g N_VDD_Mp9@2071_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2070 N_OUT9_Mp9@2070_d N_OUT8_Mp9@2070_g N_VDD_Mp9@2070_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2069 N_OUT9_Mn9@2069_d N_OUT8_Mn9@2069_g N_VSS_Mn9@2069_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2068 N_OUT9_Mn9@2068_d N_OUT8_Mn9@2068_g N_VSS_Mn9@2068_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2069 N_OUT9_Mp9@2069_d N_OUT8_Mp9@2069_g N_VDD_Mp9@2069_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2068 N_OUT9_Mp9@2068_d N_OUT8_Mp9@2068_g N_VDD_Mp9@2068_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2067 N_OUT9_Mn9@2067_d N_OUT8_Mn9@2067_g N_VSS_Mn9@2067_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2066 N_OUT9_Mn9@2066_d N_OUT8_Mn9@2066_g N_VSS_Mn9@2066_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2067 N_OUT9_Mp9@2067_d N_OUT8_Mp9@2067_g N_VDD_Mp9@2067_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2066 N_OUT9_Mp9@2066_d N_OUT8_Mp9@2066_g N_VDD_Mp9@2066_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2065 N_OUT9_Mn9@2065_d N_OUT8_Mn9@2065_g N_VSS_Mn9@2065_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2064 N_OUT9_Mn9@2064_d N_OUT8_Mn9@2064_g N_VSS_Mn9@2064_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2065 N_OUT9_Mp9@2065_d N_OUT8_Mp9@2065_g N_VDD_Mp9@2065_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2064 N_OUT9_Mp9@2064_d N_OUT8_Mp9@2064_g N_VDD_Mp9@2064_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2063 N_OUT9_Mn9@2063_d N_OUT8_Mn9@2063_g N_VSS_Mn9@2063_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2062 N_OUT9_Mn9@2062_d N_OUT8_Mn9@2062_g N_VSS_Mn9@2062_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2063 N_OUT9_Mp9@2063_d N_OUT8_Mp9@2063_g N_VDD_Mp9@2063_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2062 N_OUT9_Mp9@2062_d N_OUT8_Mp9@2062_g N_VDD_Mp9@2062_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2061 N_OUT9_Mn9@2061_d N_OUT8_Mn9@2061_g N_VSS_Mn9@2061_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2060 N_OUT9_Mn9@2060_d N_OUT8_Mn9@2060_g N_VSS_Mn9@2060_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2061 N_OUT9_Mp9@2061_d N_OUT8_Mp9@2061_g N_VDD_Mp9@2061_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2060 N_OUT9_Mp9@2060_d N_OUT8_Mp9@2060_g N_VDD_Mp9@2060_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2059 N_OUT9_Mn9@2059_d N_OUT8_Mn9@2059_g N_VSS_Mn9@2059_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2058 N_OUT9_Mn9@2058_d N_OUT8_Mn9@2058_g N_VSS_Mn9@2058_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2059 N_OUT9_Mp9@2059_d N_OUT8_Mp9@2059_g N_VDD_Mp9@2059_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2058 N_OUT9_Mp9@2058_d N_OUT8_Mp9@2058_g N_VDD_Mp9@2058_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2057 N_OUT9_Mn9@2057_d N_OUT8_Mn9@2057_g N_VSS_Mn9@2057_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2056 N_OUT9_Mn9@2056_d N_OUT8_Mn9@2056_g N_VSS_Mn9@2056_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2057 N_OUT9_Mp9@2057_d N_OUT8_Mp9@2057_g N_VDD_Mp9@2057_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2056 N_OUT9_Mp9@2056_d N_OUT8_Mp9@2056_g N_VDD_Mp9@2056_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2055 N_OUT9_Mn9@2055_d N_OUT8_Mn9@2055_g N_VSS_Mn9@2055_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2054 N_OUT9_Mn9@2054_d N_OUT8_Mn9@2054_g N_VSS_Mn9@2054_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2055 N_OUT9_Mp9@2055_d N_OUT8_Mp9@2055_g N_VDD_Mp9@2055_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2054 N_OUT9_Mp9@2054_d N_OUT8_Mp9@2054_g N_VDD_Mp9@2054_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2053 N_OUT9_Mn9@2053_d N_OUT8_Mn9@2053_g N_VSS_Mn9@2053_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2052 N_OUT9_Mn9@2052_d N_OUT8_Mn9@2052_g N_VSS_Mn9@2052_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2053 N_OUT9_Mp9@2053_d N_OUT8_Mp9@2053_g N_VDD_Mp9@2053_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2052 N_OUT9_Mp9@2052_d N_OUT8_Mp9@2052_g N_VDD_Mp9@2052_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2051 N_OUT9_Mn9@2051_d N_OUT8_Mn9@2051_g N_VSS_Mn9@2051_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2050 N_OUT9_Mn9@2050_d N_OUT8_Mn9@2050_g N_VSS_Mn9@2050_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2051 N_OUT9_Mp9@2051_d N_OUT8_Mp9@2051_g N_VDD_Mp9@2051_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2050 N_OUT9_Mp9@2050_d N_OUT8_Mp9@2050_g N_VDD_Mp9@2050_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2049 N_OUT9_Mn9@2049_d N_OUT8_Mn9@2049_g N_VSS_Mn9@2049_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2048 N_OUT9_Mn9@2048_d N_OUT8_Mn9@2048_g N_VSS_Mn9@2048_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2049 N_OUT9_Mp9@2049_d N_OUT8_Mp9@2049_g N_VDD_Mp9@2049_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2048 N_OUT9_Mp9@2048_d N_OUT8_Mp9@2048_g N_VDD_Mp9@2048_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2047 N_OUT9_Mn9@2047_d N_OUT8_Mn9@2047_g N_VSS_Mn9@2047_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2046 N_OUT9_Mn9@2046_d N_OUT8_Mn9@2046_g N_VSS_Mn9@2046_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2047 N_OUT9_Mp9@2047_d N_OUT8_Mp9@2047_g N_VDD_Mp9@2047_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2046 N_OUT9_Mp9@2046_d N_OUT8_Mp9@2046_g N_VDD_Mp9@2046_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2045 N_OUT9_Mn9@2045_d N_OUT8_Mn9@2045_g N_VSS_Mn9@2045_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2044 N_OUT9_Mn9@2044_d N_OUT8_Mn9@2044_g N_VSS_Mn9@2044_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2045 N_OUT9_Mp9@2045_d N_OUT8_Mp9@2045_g N_VDD_Mp9@2045_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2044 N_OUT9_Mp9@2044_d N_OUT8_Mp9@2044_g N_VDD_Mp9@2044_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2043 N_OUT9_Mn9@2043_d N_OUT8_Mn9@2043_g N_VSS_Mn9@2043_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2042 N_OUT9_Mn9@2042_d N_OUT8_Mn9@2042_g N_VSS_Mn9@2042_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2043 N_OUT9_Mp9@2043_d N_OUT8_Mp9@2043_g N_VDD_Mp9@2043_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2042 N_OUT9_Mp9@2042_d N_OUT8_Mp9@2042_g N_VDD_Mp9@2042_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2041 N_OUT9_Mn9@2041_d N_OUT8_Mn9@2041_g N_VSS_Mn9@2041_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2040 N_OUT9_Mn9@2040_d N_OUT8_Mn9@2040_g N_VSS_Mn9@2040_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2041 N_OUT9_Mp9@2041_d N_OUT8_Mp9@2041_g N_VDD_Mp9@2041_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2040 N_OUT9_Mp9@2040_d N_OUT8_Mp9@2040_g N_VDD_Mp9@2040_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2039 N_OUT9_Mn9@2039_d N_OUT8_Mn9@2039_g N_VSS_Mn9@2039_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2038 N_OUT9_Mn9@2038_d N_OUT8_Mn9@2038_g N_VSS_Mn9@2038_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2039 N_OUT9_Mp9@2039_d N_OUT8_Mp9@2039_g N_VDD_Mp9@2039_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2038 N_OUT9_Mp9@2038_d N_OUT8_Mp9@2038_g N_VDD_Mp9@2038_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2037 N_OUT9_Mn9@2037_d N_OUT8_Mn9@2037_g N_VSS_Mn9@2037_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2036 N_OUT9_Mn9@2036_d N_OUT8_Mn9@2036_g N_VSS_Mn9@2036_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2037 N_OUT9_Mp9@2037_d N_OUT8_Mp9@2037_g N_VDD_Mp9@2037_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2036 N_OUT9_Mp9@2036_d N_OUT8_Mp9@2036_g N_VDD_Mp9@2036_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2035 N_OUT9_Mn9@2035_d N_OUT8_Mn9@2035_g N_VSS_Mn9@2035_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2034 N_OUT9_Mn9@2034_d N_OUT8_Mn9@2034_g N_VSS_Mn9@2034_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2035 N_OUT9_Mp9@2035_d N_OUT8_Mp9@2035_g N_VDD_Mp9@2035_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2034 N_OUT9_Mp9@2034_d N_OUT8_Mp9@2034_g N_VDD_Mp9@2034_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2033 N_OUT9_Mn9@2033_d N_OUT8_Mn9@2033_g N_VSS_Mn9@2033_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2032 N_OUT9_Mn9@2032_d N_OUT8_Mn9@2032_g N_VSS_Mn9@2032_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2033 N_OUT9_Mp9@2033_d N_OUT8_Mp9@2033_g N_VDD_Mp9@2033_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2032 N_OUT9_Mp9@2032_d N_OUT8_Mp9@2032_g N_VDD_Mp9@2032_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2031 N_OUT9_Mn9@2031_d N_OUT8_Mn9@2031_g N_VSS_Mn9@2031_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2030 N_OUT9_Mn9@2030_d N_OUT8_Mn9@2030_g N_VSS_Mn9@2030_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2031 N_OUT9_Mp9@2031_d N_OUT8_Mp9@2031_g N_VDD_Mp9@2031_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2030 N_OUT9_Mp9@2030_d N_OUT8_Mp9@2030_g N_VDD_Mp9@2030_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2029 N_OUT9_Mn9@2029_d N_OUT8_Mn9@2029_g N_VSS_Mn9@2029_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2028 N_OUT9_Mn9@2028_d N_OUT8_Mn9@2028_g N_VSS_Mn9@2028_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2029 N_OUT9_Mp9@2029_d N_OUT8_Mp9@2029_g N_VDD_Mp9@2029_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2028 N_OUT9_Mp9@2028_d N_OUT8_Mp9@2028_g N_VDD_Mp9@2028_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2027 N_OUT9_Mn9@2027_d N_OUT8_Mn9@2027_g N_VSS_Mn9@2027_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2026 N_OUT9_Mn9@2026_d N_OUT8_Mn9@2026_g N_VSS_Mn9@2026_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2027 N_OUT9_Mp9@2027_d N_OUT8_Mp9@2027_g N_VDD_Mp9@2027_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2026 N_OUT9_Mp9@2026_d N_OUT8_Mp9@2026_g N_VDD_Mp9@2026_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2025 N_OUT9_Mn9@2025_d N_OUT8_Mn9@2025_g N_VSS_Mn9@2025_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2024 N_OUT9_Mn9@2024_d N_OUT8_Mn9@2024_g N_VSS_Mn9@2024_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2025 N_OUT9_Mp9@2025_d N_OUT8_Mp9@2025_g N_VDD_Mp9@2025_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2024 N_OUT9_Mp9@2024_d N_OUT8_Mp9@2024_g N_VDD_Mp9@2024_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2023 N_OUT9_Mn9@2023_d N_OUT8_Mn9@2023_g N_VSS_Mn9@2023_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2022 N_OUT9_Mn9@2022_d N_OUT8_Mn9@2022_g N_VSS_Mn9@2022_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2023 N_OUT9_Mp9@2023_d N_OUT8_Mp9@2023_g N_VDD_Mp9@2023_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2022 N_OUT9_Mp9@2022_d N_OUT8_Mp9@2022_g N_VDD_Mp9@2022_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2021 N_OUT9_Mn9@2021_d N_OUT8_Mn9@2021_g N_VSS_Mn9@2021_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2020 N_OUT9_Mn9@2020_d N_OUT8_Mn9@2020_g N_VSS_Mn9@2020_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2021 N_OUT9_Mp9@2021_d N_OUT8_Mp9@2021_g N_VDD_Mp9@2021_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2020 N_OUT9_Mp9@2020_d N_OUT8_Mp9@2020_g N_VDD_Mp9@2020_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2019 N_OUT9_Mn9@2019_d N_OUT8_Mn9@2019_g N_VSS_Mn9@2019_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2018 N_OUT9_Mn9@2018_d N_OUT8_Mn9@2018_g N_VSS_Mn9@2018_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2019 N_OUT9_Mp9@2019_d N_OUT8_Mp9@2019_g N_VDD_Mp9@2019_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2018 N_OUT9_Mp9@2018_d N_OUT8_Mp9@2018_g N_VDD_Mp9@2018_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2017 N_OUT9_Mn9@2017_d N_OUT8_Mn9@2017_g N_VSS_Mn9@2017_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2016 N_OUT9_Mn9@2016_d N_OUT8_Mn9@2016_g N_VSS_Mn9@2016_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2017 N_OUT9_Mp9@2017_d N_OUT8_Mp9@2017_g N_VDD_Mp9@2017_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2016 N_OUT9_Mp9@2016_d N_OUT8_Mp9@2016_g N_VDD_Mp9@2016_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2015 N_OUT9_Mn9@2015_d N_OUT8_Mn9@2015_g N_VSS_Mn9@2015_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2014 N_OUT9_Mn9@2014_d N_OUT8_Mn9@2014_g N_VSS_Mn9@2014_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2015 N_OUT9_Mp9@2015_d N_OUT8_Mp9@2015_g N_VDD_Mp9@2015_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2014 N_OUT9_Mp9@2014_d N_OUT8_Mp9@2014_g N_VDD_Mp9@2014_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2013 N_OUT9_Mn9@2013_d N_OUT8_Mn9@2013_g N_VSS_Mn9@2013_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2012 N_OUT9_Mn9@2012_d N_OUT8_Mn9@2012_g N_VSS_Mn9@2012_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2013 N_OUT9_Mp9@2013_d N_OUT8_Mp9@2013_g N_VDD_Mp9@2013_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2012 N_OUT9_Mp9@2012_d N_OUT8_Mp9@2012_g N_VDD_Mp9@2012_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2011 N_OUT9_Mn9@2011_d N_OUT8_Mn9@2011_g N_VSS_Mn9@2011_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2010 N_OUT9_Mn9@2010_d N_OUT8_Mn9@2010_g N_VSS_Mn9@2010_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2011 N_OUT9_Mp9@2011_d N_OUT8_Mp9@2011_g N_VDD_Mp9@2011_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2010 N_OUT9_Mp9@2010_d N_OUT8_Mp9@2010_g N_VDD_Mp9@2010_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2009 N_OUT9_Mn9@2009_d N_OUT8_Mn9@2009_g N_VSS_Mn9@2009_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2008 N_OUT9_Mn9@2008_d N_OUT8_Mn9@2008_g N_VSS_Mn9@2008_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2009 N_OUT9_Mp9@2009_d N_OUT8_Mp9@2009_g N_VDD_Mp9@2009_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2008 N_OUT9_Mp9@2008_d N_OUT8_Mp9@2008_g N_VDD_Mp9@2008_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2007 N_OUT9_Mn9@2007_d N_OUT8_Mn9@2007_g N_VSS_Mn9@2007_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2006 N_OUT9_Mn9@2006_d N_OUT8_Mn9@2006_g N_VSS_Mn9@2006_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2007 N_OUT9_Mp9@2007_d N_OUT8_Mp9@2007_g N_VDD_Mp9@2007_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2006 N_OUT9_Mp9@2006_d N_OUT8_Mp9@2006_g N_VDD_Mp9@2006_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2005 N_OUT9_Mn9@2005_d N_OUT8_Mn9@2005_g N_VSS_Mn9@2005_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2004 N_OUT9_Mn9@2004_d N_OUT8_Mn9@2004_g N_VSS_Mn9@2004_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2005 N_OUT9_Mp9@2005_d N_OUT8_Mp9@2005_g N_VDD_Mp9@2005_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2004 N_OUT9_Mp9@2004_d N_OUT8_Mp9@2004_g N_VDD_Mp9@2004_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2003 N_OUT9_Mn9@2003_d N_OUT8_Mn9@2003_g N_VSS_Mn9@2003_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2002 N_OUT9_Mn9@2002_d N_OUT8_Mn9@2002_g N_VSS_Mn9@2002_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2003 N_OUT9_Mp9@2003_d N_OUT8_Mp9@2003_g N_VDD_Mp9@2003_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2002 N_OUT9_Mp9@2002_d N_OUT8_Mp9@2002_g N_VDD_Mp9@2002_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@2001 N_OUT9_Mn9@2001_d N_OUT8_Mn9@2001_g N_VSS_Mn9@2001_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2000 N_OUT9_Mn9@2000_d N_OUT8_Mn9@2000_g N_VSS_Mn9@2000_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@2001 N_OUT9_Mp9@2001_d N_OUT8_Mp9@2001_g N_VDD_Mp9@2001_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2000 N_OUT9_Mp9@2000_d N_OUT8_Mp9@2000_g N_VDD_Mp9@2000_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1999 N_OUT9_Mn9@1999_d N_OUT8_Mn9@1999_g N_VSS_Mn9@1999_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1998 N_OUT9_Mn9@1998_d N_OUT8_Mn9@1998_g N_VSS_Mn9@1998_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1999 N_OUT9_Mp9@1999_d N_OUT8_Mp9@1999_g N_VDD_Mp9@1999_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1998 N_OUT9_Mp9@1998_d N_OUT8_Mp9@1998_g N_VDD_Mp9@1998_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1997 N_OUT9_Mn9@1997_d N_OUT8_Mn9@1997_g N_VSS_Mn9@1997_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1996 N_OUT9_Mn9@1996_d N_OUT8_Mn9@1996_g N_VSS_Mn9@1996_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1997 N_OUT9_Mp9@1997_d N_OUT8_Mp9@1997_g N_VDD_Mp9@1997_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1996 N_OUT9_Mp9@1996_d N_OUT8_Mp9@1996_g N_VDD_Mp9@1996_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1995 N_OUT9_Mn9@1995_d N_OUT8_Mn9@1995_g N_VSS_Mn9@1995_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1994 N_OUT9_Mn9@1994_d N_OUT8_Mn9@1994_g N_VSS_Mn9@1994_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1995 N_OUT9_Mp9@1995_d N_OUT8_Mp9@1995_g N_VDD_Mp9@1995_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1994 N_OUT9_Mp9@1994_d N_OUT8_Mp9@1994_g N_VDD_Mp9@1994_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1993 N_OUT9_Mn9@1993_d N_OUT8_Mn9@1993_g N_VSS_Mn9@1993_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1992 N_OUT9_Mn9@1992_d N_OUT8_Mn9@1992_g N_VSS_Mn9@1992_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1993 N_OUT9_Mp9@1993_d N_OUT8_Mp9@1993_g N_VDD_Mp9@1993_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1992 N_OUT9_Mp9@1992_d N_OUT8_Mp9@1992_g N_VDD_Mp9@1992_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1991 N_OUT9_Mn9@1991_d N_OUT8_Mn9@1991_g N_VSS_Mn9@1991_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1990 N_OUT9_Mn9@1990_d N_OUT8_Mn9@1990_g N_VSS_Mn9@1990_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1991 N_OUT9_Mp9@1991_d N_OUT8_Mp9@1991_g N_VDD_Mp9@1991_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1990 N_OUT9_Mp9@1990_d N_OUT8_Mp9@1990_g N_VDD_Mp9@1990_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1989 N_OUT9_Mn9@1989_d N_OUT8_Mn9@1989_g N_VSS_Mn9@1989_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1988 N_OUT9_Mn9@1988_d N_OUT8_Mn9@1988_g N_VSS_Mn9@1988_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1989 N_OUT9_Mp9@1989_d N_OUT8_Mp9@1989_g N_VDD_Mp9@1989_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1988 N_OUT9_Mp9@1988_d N_OUT8_Mp9@1988_g N_VDD_Mp9@1988_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1987 N_OUT9_Mn9@1987_d N_OUT8_Mn9@1987_g N_VSS_Mn9@1987_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1986 N_OUT9_Mn9@1986_d N_OUT8_Mn9@1986_g N_VSS_Mn9@1986_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1987 N_OUT9_Mp9@1987_d N_OUT8_Mp9@1987_g N_VDD_Mp9@1987_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1986 N_OUT9_Mp9@1986_d N_OUT8_Mp9@1986_g N_VDD_Mp9@1986_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1985 N_OUT9_Mn9@1985_d N_OUT8_Mn9@1985_g N_VSS_Mn9@1985_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1984 N_OUT9_Mn9@1984_d N_OUT8_Mn9@1984_g N_VSS_Mn9@1984_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1985 N_OUT9_Mp9@1985_d N_OUT8_Mp9@1985_g N_VDD_Mp9@1985_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1984 N_OUT9_Mp9@1984_d N_OUT8_Mp9@1984_g N_VDD_Mp9@1984_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1983 N_OUT9_Mn9@1983_d N_OUT8_Mn9@1983_g N_VSS_Mn9@1983_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1982 N_OUT9_Mn9@1982_d N_OUT8_Mn9@1982_g N_VSS_Mn9@1982_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1983 N_OUT9_Mp9@1983_d N_OUT8_Mp9@1983_g N_VDD_Mp9@1983_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1982 N_OUT9_Mp9@1982_d N_OUT8_Mp9@1982_g N_VDD_Mp9@1982_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1981 N_OUT9_Mn9@1981_d N_OUT8_Mn9@1981_g N_VSS_Mn9@1981_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1980 N_OUT9_Mn9@1980_d N_OUT8_Mn9@1980_g N_VSS_Mn9@1980_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1981 N_OUT9_Mp9@1981_d N_OUT8_Mp9@1981_g N_VDD_Mp9@1981_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1980 N_OUT9_Mp9@1980_d N_OUT8_Mp9@1980_g N_VDD_Mp9@1980_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1979 N_OUT9_Mn9@1979_d N_OUT8_Mn9@1979_g N_VSS_Mn9@1979_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1978 N_OUT9_Mn9@1978_d N_OUT8_Mn9@1978_g N_VSS_Mn9@1978_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1979 N_OUT9_Mp9@1979_d N_OUT8_Mp9@1979_g N_VDD_Mp9@1979_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1978 N_OUT9_Mp9@1978_d N_OUT8_Mp9@1978_g N_VDD_Mp9@1978_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1977 N_OUT9_Mn9@1977_d N_OUT8_Mn9@1977_g N_VSS_Mn9@1977_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1976 N_OUT9_Mn9@1976_d N_OUT8_Mn9@1976_g N_VSS_Mn9@1976_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1977 N_OUT9_Mp9@1977_d N_OUT8_Mp9@1977_g N_VDD_Mp9@1977_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1976 N_OUT9_Mp9@1976_d N_OUT8_Mp9@1976_g N_VDD_Mp9@1976_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1975 N_OUT9_Mn9@1975_d N_OUT8_Mn9@1975_g N_VSS_Mn9@1975_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1974 N_OUT9_Mn9@1974_d N_OUT8_Mn9@1974_g N_VSS_Mn9@1974_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1975 N_OUT9_Mp9@1975_d N_OUT8_Mp9@1975_g N_VDD_Mp9@1975_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1974 N_OUT9_Mp9@1974_d N_OUT8_Mp9@1974_g N_VDD_Mp9@1974_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1973 N_OUT9_Mn9@1973_d N_OUT8_Mn9@1973_g N_VSS_Mn9@1973_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1972 N_OUT9_Mn9@1972_d N_OUT8_Mn9@1972_g N_VSS_Mn9@1972_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1973 N_OUT9_Mp9@1973_d N_OUT8_Mp9@1973_g N_VDD_Mp9@1973_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1972 N_OUT9_Mp9@1972_d N_OUT8_Mp9@1972_g N_VDD_Mp9@1972_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1971 N_OUT9_Mn9@1971_d N_OUT8_Mn9@1971_g N_VSS_Mn9@1971_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1970 N_OUT9_Mn9@1970_d N_OUT8_Mn9@1970_g N_VSS_Mn9@1970_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1971 N_OUT9_Mp9@1971_d N_OUT8_Mp9@1971_g N_VDD_Mp9@1971_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1970 N_OUT9_Mp9@1970_d N_OUT8_Mp9@1970_g N_VDD_Mp9@1970_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1969 N_OUT9_Mn9@1969_d N_OUT8_Mn9@1969_g N_VSS_Mn9@1969_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1968 N_OUT9_Mn9@1968_d N_OUT8_Mn9@1968_g N_VSS_Mn9@1968_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1969 N_OUT9_Mp9@1969_d N_OUT8_Mp9@1969_g N_VDD_Mp9@1969_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1968 N_OUT9_Mp9@1968_d N_OUT8_Mp9@1968_g N_VDD_Mp9@1968_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1967 N_OUT9_Mn9@1967_d N_OUT8_Mn9@1967_g N_VSS_Mn9@1967_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1966 N_OUT9_Mn9@1966_d N_OUT8_Mn9@1966_g N_VSS_Mn9@1966_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1967 N_OUT9_Mp9@1967_d N_OUT8_Mp9@1967_g N_VDD_Mp9@1967_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1966 N_OUT9_Mp9@1966_d N_OUT8_Mp9@1966_g N_VDD_Mp9@1966_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1965 N_OUT9_Mn9@1965_d N_OUT8_Mn9@1965_g N_VSS_Mn9@1965_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1964 N_OUT9_Mn9@1964_d N_OUT8_Mn9@1964_g N_VSS_Mn9@1964_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1965 N_OUT9_Mp9@1965_d N_OUT8_Mp9@1965_g N_VDD_Mp9@1965_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1964 N_OUT9_Mp9@1964_d N_OUT8_Mp9@1964_g N_VDD_Mp9@1964_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1963 N_OUT9_Mn9@1963_d N_OUT8_Mn9@1963_g N_VSS_Mn9@1963_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1962 N_OUT9_Mn9@1962_d N_OUT8_Mn9@1962_g N_VSS_Mn9@1962_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1963 N_OUT9_Mp9@1963_d N_OUT8_Mp9@1963_g N_VDD_Mp9@1963_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1962 N_OUT9_Mp9@1962_d N_OUT8_Mp9@1962_g N_VDD_Mp9@1962_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1961 N_OUT9_Mn9@1961_d N_OUT8_Mn9@1961_g N_VSS_Mn9@1961_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1960 N_OUT9_Mn9@1960_d N_OUT8_Mn9@1960_g N_VSS_Mn9@1960_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1961 N_OUT9_Mp9@1961_d N_OUT8_Mp9@1961_g N_VDD_Mp9@1961_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1960 N_OUT9_Mp9@1960_d N_OUT8_Mp9@1960_g N_VDD_Mp9@1960_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1959 N_OUT9_Mn9@1959_d N_OUT8_Mn9@1959_g N_VSS_Mn9@1959_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1958 N_OUT9_Mn9@1958_d N_OUT8_Mn9@1958_g N_VSS_Mn9@1958_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1959 N_OUT9_Mp9@1959_d N_OUT8_Mp9@1959_g N_VDD_Mp9@1959_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1958 N_OUT9_Mp9@1958_d N_OUT8_Mp9@1958_g N_VDD_Mp9@1958_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1957 N_OUT9_Mn9@1957_d N_OUT8_Mn9@1957_g N_VSS_Mn9@1957_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1956 N_OUT9_Mn9@1956_d N_OUT8_Mn9@1956_g N_VSS_Mn9@1956_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1957 N_OUT9_Mp9@1957_d N_OUT8_Mp9@1957_g N_VDD_Mp9@1957_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1956 N_OUT9_Mp9@1956_d N_OUT8_Mp9@1956_g N_VDD_Mp9@1956_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1955 N_OUT9_Mn9@1955_d N_OUT8_Mn9@1955_g N_VSS_Mn9@1955_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1954 N_OUT9_Mn9@1954_d N_OUT8_Mn9@1954_g N_VSS_Mn9@1954_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1955 N_OUT9_Mp9@1955_d N_OUT8_Mp9@1955_g N_VDD_Mp9@1955_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1954 N_OUT9_Mp9@1954_d N_OUT8_Mp9@1954_g N_VDD_Mp9@1954_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1953 N_OUT9_Mn9@1953_d N_OUT8_Mn9@1953_g N_VSS_Mn9@1953_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1952 N_OUT9_Mn9@1952_d N_OUT8_Mn9@1952_g N_VSS_Mn9@1952_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1953 N_OUT9_Mp9@1953_d N_OUT8_Mp9@1953_g N_VDD_Mp9@1953_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1952 N_OUT9_Mp9@1952_d N_OUT8_Mp9@1952_g N_VDD_Mp9@1952_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1951 N_OUT9_Mn9@1951_d N_OUT8_Mn9@1951_g N_VSS_Mn9@1951_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1950 N_OUT9_Mn9@1950_d N_OUT8_Mn9@1950_g N_VSS_Mn9@1950_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1951 N_OUT9_Mp9@1951_d N_OUT8_Mp9@1951_g N_VDD_Mp9@1951_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1950 N_OUT9_Mp9@1950_d N_OUT8_Mp9@1950_g N_VDD_Mp9@1950_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1949 N_OUT9_Mn9@1949_d N_OUT8_Mn9@1949_g N_VSS_Mn9@1949_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1948 N_OUT9_Mn9@1948_d N_OUT8_Mn9@1948_g N_VSS_Mn9@1948_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1949 N_OUT9_Mp9@1949_d N_OUT8_Mp9@1949_g N_VDD_Mp9@1949_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1948 N_OUT9_Mp9@1948_d N_OUT8_Mp9@1948_g N_VDD_Mp9@1948_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1947 N_OUT9_Mn9@1947_d N_OUT8_Mn9@1947_g N_VSS_Mn9@1947_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1946 N_OUT9_Mn9@1946_d N_OUT8_Mn9@1946_g N_VSS_Mn9@1946_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1947 N_OUT9_Mp9@1947_d N_OUT8_Mp9@1947_g N_VDD_Mp9@1947_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1946 N_OUT9_Mp9@1946_d N_OUT8_Mp9@1946_g N_VDD_Mp9@1946_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1945 N_OUT9_Mn9@1945_d N_OUT8_Mn9@1945_g N_VSS_Mn9@1945_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1944 N_OUT9_Mn9@1944_d N_OUT8_Mn9@1944_g N_VSS_Mn9@1944_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1945 N_OUT9_Mp9@1945_d N_OUT8_Mp9@1945_g N_VDD_Mp9@1945_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1944 N_OUT9_Mp9@1944_d N_OUT8_Mp9@1944_g N_VDD_Mp9@1944_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1943 N_OUT9_Mn9@1943_d N_OUT8_Mn9@1943_g N_VSS_Mn9@1943_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1942 N_OUT9_Mn9@1942_d N_OUT8_Mn9@1942_g N_VSS_Mn9@1942_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1943 N_OUT9_Mp9@1943_d N_OUT8_Mp9@1943_g N_VDD_Mp9@1943_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1942 N_OUT9_Mp9@1942_d N_OUT8_Mp9@1942_g N_VDD_Mp9@1942_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1941 N_OUT9_Mn9@1941_d N_OUT8_Mn9@1941_g N_VSS_Mn9@1941_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1940 N_OUT9_Mn9@1940_d N_OUT8_Mn9@1940_g N_VSS_Mn9@1940_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1941 N_OUT9_Mp9@1941_d N_OUT8_Mp9@1941_g N_VDD_Mp9@1941_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1940 N_OUT9_Mp9@1940_d N_OUT8_Mp9@1940_g N_VDD_Mp9@1940_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1939 N_OUT9_Mn9@1939_d N_OUT8_Mn9@1939_g N_VSS_Mn9@1939_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1938 N_OUT9_Mn9@1938_d N_OUT8_Mn9@1938_g N_VSS_Mn9@1938_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1939 N_OUT9_Mp9@1939_d N_OUT8_Mp9@1939_g N_VDD_Mp9@1939_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1938 N_OUT9_Mp9@1938_d N_OUT8_Mp9@1938_g N_VDD_Mp9@1938_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1937 N_OUT9_Mn9@1937_d N_OUT8_Mn9@1937_g N_VSS_Mn9@1937_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1936 N_OUT9_Mn9@1936_d N_OUT8_Mn9@1936_g N_VSS_Mn9@1936_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1937 N_OUT9_Mp9@1937_d N_OUT8_Mp9@1937_g N_VDD_Mp9@1937_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1936 N_OUT9_Mp9@1936_d N_OUT8_Mp9@1936_g N_VDD_Mp9@1936_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1935 N_OUT9_Mn9@1935_d N_OUT8_Mn9@1935_g N_VSS_Mn9@1935_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1934 N_OUT9_Mn9@1934_d N_OUT8_Mn9@1934_g N_VSS_Mn9@1934_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1935 N_OUT9_Mp9@1935_d N_OUT8_Mp9@1935_g N_VDD_Mp9@1935_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1934 N_OUT9_Mp9@1934_d N_OUT8_Mp9@1934_g N_VDD_Mp9@1934_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1933 N_OUT9_Mn9@1933_d N_OUT8_Mn9@1933_g N_VSS_Mn9@1933_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1932 N_OUT9_Mn9@1932_d N_OUT8_Mn9@1932_g N_VSS_Mn9@1932_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1933 N_OUT9_Mp9@1933_d N_OUT8_Mp9@1933_g N_VDD_Mp9@1933_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1932 N_OUT9_Mp9@1932_d N_OUT8_Mp9@1932_g N_VDD_Mp9@1932_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1931 N_OUT9_Mn9@1931_d N_OUT8_Mn9@1931_g N_VSS_Mn9@1931_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1930 N_OUT9_Mn9@1930_d N_OUT8_Mn9@1930_g N_VSS_Mn9@1930_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1931 N_OUT9_Mp9@1931_d N_OUT8_Mp9@1931_g N_VDD_Mp9@1931_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1930 N_OUT9_Mp9@1930_d N_OUT8_Mp9@1930_g N_VDD_Mp9@1930_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1929 N_OUT9_Mn9@1929_d N_OUT8_Mn9@1929_g N_VSS_Mn9@1929_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1928 N_OUT9_Mn9@1928_d N_OUT8_Mn9@1928_g N_VSS_Mn9@1928_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1929 N_OUT9_Mp9@1929_d N_OUT8_Mp9@1929_g N_VDD_Mp9@1929_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1928 N_OUT9_Mp9@1928_d N_OUT8_Mp9@1928_g N_VDD_Mp9@1928_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1927 N_OUT9_Mn9@1927_d N_OUT8_Mn9@1927_g N_VSS_Mn9@1927_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1926 N_OUT9_Mn9@1926_d N_OUT8_Mn9@1926_g N_VSS_Mn9@1926_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1927 N_OUT9_Mp9@1927_d N_OUT8_Mp9@1927_g N_VDD_Mp9@1927_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1926 N_OUT9_Mp9@1926_d N_OUT8_Mp9@1926_g N_VDD_Mp9@1926_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1925 N_OUT9_Mn9@1925_d N_OUT8_Mn9@1925_g N_VSS_Mn9@1925_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1924 N_OUT9_Mn9@1924_d N_OUT8_Mn9@1924_g N_VSS_Mn9@1924_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1925 N_OUT9_Mp9@1925_d N_OUT8_Mp9@1925_g N_VDD_Mp9@1925_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1924 N_OUT9_Mp9@1924_d N_OUT8_Mp9@1924_g N_VDD_Mp9@1924_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1923 N_OUT9_Mn9@1923_d N_OUT8_Mn9@1923_g N_VSS_Mn9@1923_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1922 N_OUT9_Mn9@1922_d N_OUT8_Mn9@1922_g N_VSS_Mn9@1922_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1923 N_OUT9_Mp9@1923_d N_OUT8_Mp9@1923_g N_VDD_Mp9@1923_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1922 N_OUT9_Mp9@1922_d N_OUT8_Mp9@1922_g N_VDD_Mp9@1922_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1921 N_OUT9_Mn9@1921_d N_OUT8_Mn9@1921_g N_VSS_Mn9@1921_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1920 N_OUT9_Mn9@1920_d N_OUT8_Mn9@1920_g N_VSS_Mn9@1920_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1921 N_OUT9_Mp9@1921_d N_OUT8_Mp9@1921_g N_VDD_Mp9@1921_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1920 N_OUT9_Mp9@1920_d N_OUT8_Mp9@1920_g N_VDD_Mp9@1920_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1919 N_OUT9_Mn9@1919_d N_OUT8_Mn9@1919_g N_VSS_Mn9@1919_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1918 N_OUT9_Mn9@1918_d N_OUT8_Mn9@1918_g N_VSS_Mn9@1918_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1919 N_OUT9_Mp9@1919_d N_OUT8_Mp9@1919_g N_VDD_Mp9@1919_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1918 N_OUT9_Mp9@1918_d N_OUT8_Mp9@1918_g N_VDD_Mp9@1918_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1917 N_OUT9_Mn9@1917_d N_OUT8_Mn9@1917_g N_VSS_Mn9@1917_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1916 N_OUT9_Mn9@1916_d N_OUT8_Mn9@1916_g N_VSS_Mn9@1916_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1917 N_OUT9_Mp9@1917_d N_OUT8_Mp9@1917_g N_VDD_Mp9@1917_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1916 N_OUT9_Mp9@1916_d N_OUT8_Mp9@1916_g N_VDD_Mp9@1916_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1915 N_OUT9_Mn9@1915_d N_OUT8_Mn9@1915_g N_VSS_Mn9@1915_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1914 N_OUT9_Mn9@1914_d N_OUT8_Mn9@1914_g N_VSS_Mn9@1914_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1915 N_OUT9_Mp9@1915_d N_OUT8_Mp9@1915_g N_VDD_Mp9@1915_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1914 N_OUT9_Mp9@1914_d N_OUT8_Mp9@1914_g N_VDD_Mp9@1914_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1913 N_OUT9_Mn9@1913_d N_OUT8_Mn9@1913_g N_VSS_Mn9@1913_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1912 N_OUT9_Mn9@1912_d N_OUT8_Mn9@1912_g N_VSS_Mn9@1912_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1913 N_OUT9_Mp9@1913_d N_OUT8_Mp9@1913_g N_VDD_Mp9@1913_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1912 N_OUT9_Mp9@1912_d N_OUT8_Mp9@1912_g N_VDD_Mp9@1912_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1911 N_OUT9_Mn9@1911_d N_OUT8_Mn9@1911_g N_VSS_Mn9@1911_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1910 N_OUT9_Mn9@1910_d N_OUT8_Mn9@1910_g N_VSS_Mn9@1910_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1911 N_OUT9_Mp9@1911_d N_OUT8_Mp9@1911_g N_VDD_Mp9@1911_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1910 N_OUT9_Mp9@1910_d N_OUT8_Mp9@1910_g N_VDD_Mp9@1910_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1909 N_OUT9_Mn9@1909_d N_OUT8_Mn9@1909_g N_VSS_Mn9@1909_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1908 N_OUT9_Mn9@1908_d N_OUT8_Mn9@1908_g N_VSS_Mn9@1908_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1909 N_OUT9_Mp9@1909_d N_OUT8_Mp9@1909_g N_VDD_Mp9@1909_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1908 N_OUT9_Mp9@1908_d N_OUT8_Mp9@1908_g N_VDD_Mp9@1908_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1907 N_OUT9_Mn9@1907_d N_OUT8_Mn9@1907_g N_VSS_Mn9@1907_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1906 N_OUT9_Mn9@1906_d N_OUT8_Mn9@1906_g N_VSS_Mn9@1906_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1907 N_OUT9_Mp9@1907_d N_OUT8_Mp9@1907_g N_VDD_Mp9@1907_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1906 N_OUT9_Mp9@1906_d N_OUT8_Mp9@1906_g N_VDD_Mp9@1906_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1905 N_OUT9_Mn9@1905_d N_OUT8_Mn9@1905_g N_VSS_Mn9@1905_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1904 N_OUT9_Mn9@1904_d N_OUT8_Mn9@1904_g N_VSS_Mn9@1904_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1905 N_OUT9_Mp9@1905_d N_OUT8_Mp9@1905_g N_VDD_Mp9@1905_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1904 N_OUT9_Mp9@1904_d N_OUT8_Mp9@1904_g N_VDD_Mp9@1904_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1903 N_OUT9_Mn9@1903_d N_OUT8_Mn9@1903_g N_VSS_Mn9@1903_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1902 N_OUT9_Mn9@1902_d N_OUT8_Mn9@1902_g N_VSS_Mn9@1902_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1903 N_OUT9_Mp9@1903_d N_OUT8_Mp9@1903_g N_VDD_Mp9@1903_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1902 N_OUT9_Mp9@1902_d N_OUT8_Mp9@1902_g N_VDD_Mp9@1902_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1901 N_OUT9_Mn9@1901_d N_OUT8_Mn9@1901_g N_VSS_Mn9@1901_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1900 N_OUT9_Mn9@1900_d N_OUT8_Mn9@1900_g N_VSS_Mn9@1900_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1901 N_OUT9_Mp9@1901_d N_OUT8_Mp9@1901_g N_VDD_Mp9@1901_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1900 N_OUT9_Mp9@1900_d N_OUT8_Mp9@1900_g N_VDD_Mp9@1900_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1899 N_OUT9_Mn9@1899_d N_OUT8_Mn9@1899_g N_VSS_Mn9@1899_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1898 N_OUT9_Mn9@1898_d N_OUT8_Mn9@1898_g N_VSS_Mn9@1898_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1899 N_OUT9_Mp9@1899_d N_OUT8_Mp9@1899_g N_VDD_Mp9@1899_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1898 N_OUT9_Mp9@1898_d N_OUT8_Mp9@1898_g N_VDD_Mp9@1898_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1897 N_OUT9_Mn9@1897_d N_OUT8_Mn9@1897_g N_VSS_Mn9@1897_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1896 N_OUT9_Mn9@1896_d N_OUT8_Mn9@1896_g N_VSS_Mn9@1896_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1897 N_OUT9_Mp9@1897_d N_OUT8_Mp9@1897_g N_VDD_Mp9@1897_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1896 N_OUT9_Mp9@1896_d N_OUT8_Mp9@1896_g N_VDD_Mp9@1896_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1895 N_OUT9_Mn9@1895_d N_OUT8_Mn9@1895_g N_VSS_Mn9@1895_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1894 N_OUT9_Mn9@1894_d N_OUT8_Mn9@1894_g N_VSS_Mn9@1894_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1895 N_OUT9_Mp9@1895_d N_OUT8_Mp9@1895_g N_VDD_Mp9@1895_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1894 N_OUT9_Mp9@1894_d N_OUT8_Mp9@1894_g N_VDD_Mp9@1894_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1893 N_OUT9_Mn9@1893_d N_OUT8_Mn9@1893_g N_VSS_Mn9@1893_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1892 N_OUT9_Mn9@1892_d N_OUT8_Mn9@1892_g N_VSS_Mn9@1892_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1893 N_OUT9_Mp9@1893_d N_OUT8_Mp9@1893_g N_VDD_Mp9@1893_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1892 N_OUT9_Mp9@1892_d N_OUT8_Mp9@1892_g N_VDD_Mp9@1892_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1891 N_OUT9_Mn9@1891_d N_OUT8_Mn9@1891_g N_VSS_Mn9@1891_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1890 N_OUT9_Mn9@1890_d N_OUT8_Mn9@1890_g N_VSS_Mn9@1890_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1891 N_OUT9_Mp9@1891_d N_OUT8_Mp9@1891_g N_VDD_Mp9@1891_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1890 N_OUT9_Mp9@1890_d N_OUT8_Mp9@1890_g N_VDD_Mp9@1890_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1889 N_OUT9_Mn9@1889_d N_OUT8_Mn9@1889_g N_VSS_Mn9@1889_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1888 N_OUT9_Mn9@1888_d N_OUT8_Mn9@1888_g N_VSS_Mn9@1888_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1889 N_OUT9_Mp9@1889_d N_OUT8_Mp9@1889_g N_VDD_Mp9@1889_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1888 N_OUT9_Mp9@1888_d N_OUT8_Mp9@1888_g N_VDD_Mp9@1888_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1887 N_OUT9_Mn9@1887_d N_OUT8_Mn9@1887_g N_VSS_Mn9@1887_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1886 N_OUT9_Mn9@1886_d N_OUT8_Mn9@1886_g N_VSS_Mn9@1886_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1887 N_OUT9_Mp9@1887_d N_OUT8_Mp9@1887_g N_VDD_Mp9@1887_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1886 N_OUT9_Mp9@1886_d N_OUT8_Mp9@1886_g N_VDD_Mp9@1886_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1885 N_OUT9_Mn9@1885_d N_OUT8_Mn9@1885_g N_VSS_Mn9@1885_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1884 N_OUT9_Mn9@1884_d N_OUT8_Mn9@1884_g N_VSS_Mn9@1884_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1885 N_OUT9_Mp9@1885_d N_OUT8_Mp9@1885_g N_VDD_Mp9@1885_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1884 N_OUT9_Mp9@1884_d N_OUT8_Mp9@1884_g N_VDD_Mp9@1884_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1883 N_OUT9_Mn9@1883_d N_OUT8_Mn9@1883_g N_VSS_Mn9@1883_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1882 N_OUT9_Mn9@1882_d N_OUT8_Mn9@1882_g N_VSS_Mn9@1882_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1883 N_OUT9_Mp9@1883_d N_OUT8_Mp9@1883_g N_VDD_Mp9@1883_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1882 N_OUT9_Mp9@1882_d N_OUT8_Mp9@1882_g N_VDD_Mp9@1882_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1881 N_OUT9_Mn9@1881_d N_OUT8_Mn9@1881_g N_VSS_Mn9@1881_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1880 N_OUT9_Mn9@1880_d N_OUT8_Mn9@1880_g N_VSS_Mn9@1880_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1881 N_OUT9_Mp9@1881_d N_OUT8_Mp9@1881_g N_VDD_Mp9@1881_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1880 N_OUT9_Mp9@1880_d N_OUT8_Mp9@1880_g N_VDD_Mp9@1880_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1879 N_OUT9_Mn9@1879_d N_OUT8_Mn9@1879_g N_VSS_Mn9@1879_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1878 N_OUT9_Mn9@1878_d N_OUT8_Mn9@1878_g N_VSS_Mn9@1878_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1879 N_OUT9_Mp9@1879_d N_OUT8_Mp9@1879_g N_VDD_Mp9@1879_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1878 N_OUT9_Mp9@1878_d N_OUT8_Mp9@1878_g N_VDD_Mp9@1878_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1877 N_OUT9_Mn9@1877_d N_OUT8_Mn9@1877_g N_VSS_Mn9@1877_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1876 N_OUT9_Mn9@1876_d N_OUT8_Mn9@1876_g N_VSS_Mn9@1876_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1877 N_OUT9_Mp9@1877_d N_OUT8_Mp9@1877_g N_VDD_Mp9@1877_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1876 N_OUT9_Mp9@1876_d N_OUT8_Mp9@1876_g N_VDD_Mp9@1876_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1875 N_OUT9_Mn9@1875_d N_OUT8_Mn9@1875_g N_VSS_Mn9@1875_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1874 N_OUT9_Mn9@1874_d N_OUT8_Mn9@1874_g N_VSS_Mn9@1874_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1875 N_OUT9_Mp9@1875_d N_OUT8_Mp9@1875_g N_VDD_Mp9@1875_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1874 N_OUT9_Mp9@1874_d N_OUT8_Mp9@1874_g N_VDD_Mp9@1874_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1873 N_OUT9_Mn9@1873_d N_OUT8_Mn9@1873_g N_VSS_Mn9@1873_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1872 N_OUT9_Mn9@1872_d N_OUT8_Mn9@1872_g N_VSS_Mn9@1872_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1873 N_OUT9_Mp9@1873_d N_OUT8_Mp9@1873_g N_VDD_Mp9@1873_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1872 N_OUT9_Mp9@1872_d N_OUT8_Mp9@1872_g N_VDD_Mp9@1872_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1871 N_OUT9_Mn9@1871_d N_OUT8_Mn9@1871_g N_VSS_Mn9@1871_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1870 N_OUT9_Mn9@1870_d N_OUT8_Mn9@1870_g N_VSS_Mn9@1870_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1871 N_OUT9_Mp9@1871_d N_OUT8_Mp9@1871_g N_VDD_Mp9@1871_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1870 N_OUT9_Mp9@1870_d N_OUT8_Mp9@1870_g N_VDD_Mp9@1870_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1869 N_OUT9_Mn9@1869_d N_OUT8_Mn9@1869_g N_VSS_Mn9@1869_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1868 N_OUT9_Mn9@1868_d N_OUT8_Mn9@1868_g N_VSS_Mn9@1868_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1869 N_OUT9_Mp9@1869_d N_OUT8_Mp9@1869_g N_VDD_Mp9@1869_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1868 N_OUT9_Mp9@1868_d N_OUT8_Mp9@1868_g N_VDD_Mp9@1868_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1867 N_OUT9_Mn9@1867_d N_OUT8_Mn9@1867_g N_VSS_Mn9@1867_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1866 N_OUT9_Mn9@1866_d N_OUT8_Mn9@1866_g N_VSS_Mn9@1866_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1867 N_OUT9_Mp9@1867_d N_OUT8_Mp9@1867_g N_VDD_Mp9@1867_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1866 N_OUT9_Mp9@1866_d N_OUT8_Mp9@1866_g N_VDD_Mp9@1866_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1865 N_OUT9_Mn9@1865_d N_OUT8_Mn9@1865_g N_VSS_Mn9@1865_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1864 N_OUT9_Mn9@1864_d N_OUT8_Mn9@1864_g N_VSS_Mn9@1864_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1865 N_OUT9_Mp9@1865_d N_OUT8_Mp9@1865_g N_VDD_Mp9@1865_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1864 N_OUT9_Mp9@1864_d N_OUT8_Mp9@1864_g N_VDD_Mp9@1864_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1863 N_OUT9_Mn9@1863_d N_OUT8_Mn9@1863_g N_VSS_Mn9@1863_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1862 N_OUT9_Mn9@1862_d N_OUT8_Mn9@1862_g N_VSS_Mn9@1862_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1863 N_OUT9_Mp9@1863_d N_OUT8_Mp9@1863_g N_VDD_Mp9@1863_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1862 N_OUT9_Mp9@1862_d N_OUT8_Mp9@1862_g N_VDD_Mp9@1862_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1861 N_OUT9_Mn9@1861_d N_OUT8_Mn9@1861_g N_VSS_Mn9@1861_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1860 N_OUT9_Mn9@1860_d N_OUT8_Mn9@1860_g N_VSS_Mn9@1860_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1861 N_OUT9_Mp9@1861_d N_OUT8_Mp9@1861_g N_VDD_Mp9@1861_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1860 N_OUT9_Mp9@1860_d N_OUT8_Mp9@1860_g N_VDD_Mp9@1860_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1859 N_OUT9_Mn9@1859_d N_OUT8_Mn9@1859_g N_VSS_Mn9@1859_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1858 N_OUT9_Mn9@1858_d N_OUT8_Mn9@1858_g N_VSS_Mn9@1858_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1859 N_OUT9_Mp9@1859_d N_OUT8_Mp9@1859_g N_VDD_Mp9@1859_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1858 N_OUT9_Mp9@1858_d N_OUT8_Mp9@1858_g N_VDD_Mp9@1858_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1857 N_OUT9_Mn9@1857_d N_OUT8_Mn9@1857_g N_VSS_Mn9@1857_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1856 N_OUT9_Mn9@1856_d N_OUT8_Mn9@1856_g N_VSS_Mn9@1856_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1857 N_OUT9_Mp9@1857_d N_OUT8_Mp9@1857_g N_VDD_Mp9@1857_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1856 N_OUT9_Mp9@1856_d N_OUT8_Mp9@1856_g N_VDD_Mp9@1856_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1855 N_OUT9_Mn9@1855_d N_OUT8_Mn9@1855_g N_VSS_Mn9@1855_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1854 N_OUT9_Mn9@1854_d N_OUT8_Mn9@1854_g N_VSS_Mn9@1854_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1855 N_OUT9_Mp9@1855_d N_OUT8_Mp9@1855_g N_VDD_Mp9@1855_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1854 N_OUT9_Mp9@1854_d N_OUT8_Mp9@1854_g N_VDD_Mp9@1854_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1853 N_OUT9_Mn9@1853_d N_OUT8_Mn9@1853_g N_VSS_Mn9@1853_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1852 N_OUT9_Mn9@1852_d N_OUT8_Mn9@1852_g N_VSS_Mn9@1852_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1853 N_OUT9_Mp9@1853_d N_OUT8_Mp9@1853_g N_VDD_Mp9@1853_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1852 N_OUT9_Mp9@1852_d N_OUT8_Mp9@1852_g N_VDD_Mp9@1852_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1851 N_OUT9_Mn9@1851_d N_OUT8_Mn9@1851_g N_VSS_Mn9@1851_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1850 N_OUT9_Mn9@1850_d N_OUT8_Mn9@1850_g N_VSS_Mn9@1850_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1851 N_OUT9_Mp9@1851_d N_OUT8_Mp9@1851_g N_VDD_Mp9@1851_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1850 N_OUT9_Mp9@1850_d N_OUT8_Mp9@1850_g N_VDD_Mp9@1850_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1849 N_OUT9_Mn9@1849_d N_OUT8_Mn9@1849_g N_VSS_Mn9@1849_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1848 N_OUT9_Mn9@1848_d N_OUT8_Mn9@1848_g N_VSS_Mn9@1848_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1849 N_OUT9_Mp9@1849_d N_OUT8_Mp9@1849_g N_VDD_Mp9@1849_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1848 N_OUT9_Mp9@1848_d N_OUT8_Mp9@1848_g N_VDD_Mp9@1848_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1847 N_OUT9_Mn9@1847_d N_OUT8_Mn9@1847_g N_VSS_Mn9@1847_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1846 N_OUT9_Mn9@1846_d N_OUT8_Mn9@1846_g N_VSS_Mn9@1846_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1847 N_OUT9_Mp9@1847_d N_OUT8_Mp9@1847_g N_VDD_Mp9@1847_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1846 N_OUT9_Mp9@1846_d N_OUT8_Mp9@1846_g N_VDD_Mp9@1846_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1845 N_OUT9_Mn9@1845_d N_OUT8_Mn9@1845_g N_VSS_Mn9@1845_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1844 N_OUT9_Mn9@1844_d N_OUT8_Mn9@1844_g N_VSS_Mn9@1844_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1845 N_OUT9_Mp9@1845_d N_OUT8_Mp9@1845_g N_VDD_Mp9@1845_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1844 N_OUT9_Mp9@1844_d N_OUT8_Mp9@1844_g N_VDD_Mp9@1844_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1843 N_OUT9_Mn9@1843_d N_OUT8_Mn9@1843_g N_VSS_Mn9@1843_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1842 N_OUT9_Mn9@1842_d N_OUT8_Mn9@1842_g N_VSS_Mn9@1842_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1843 N_OUT9_Mp9@1843_d N_OUT8_Mp9@1843_g N_VDD_Mp9@1843_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1842 N_OUT9_Mp9@1842_d N_OUT8_Mp9@1842_g N_VDD_Mp9@1842_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1841 N_OUT9_Mn9@1841_d N_OUT8_Mn9@1841_g N_VSS_Mn9@1841_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1840 N_OUT9_Mn9@1840_d N_OUT8_Mn9@1840_g N_VSS_Mn9@1840_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1841 N_OUT9_Mp9@1841_d N_OUT8_Mp9@1841_g N_VDD_Mp9@1841_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1840 N_OUT9_Mp9@1840_d N_OUT8_Mp9@1840_g N_VDD_Mp9@1840_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1839 N_OUT9_Mn9@1839_d N_OUT8_Mn9@1839_g N_VSS_Mn9@1839_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1838 N_OUT9_Mn9@1838_d N_OUT8_Mn9@1838_g N_VSS_Mn9@1838_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1839 N_OUT9_Mp9@1839_d N_OUT8_Mp9@1839_g N_VDD_Mp9@1839_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1838 N_OUT9_Mp9@1838_d N_OUT8_Mp9@1838_g N_VDD_Mp9@1838_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1837 N_OUT9_Mn9@1837_d N_OUT8_Mn9@1837_g N_VSS_Mn9@1837_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1836 N_OUT9_Mn9@1836_d N_OUT8_Mn9@1836_g N_VSS_Mn9@1836_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1837 N_OUT9_Mp9@1837_d N_OUT8_Mp9@1837_g N_VDD_Mp9@1837_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1836 N_OUT9_Mp9@1836_d N_OUT8_Mp9@1836_g N_VDD_Mp9@1836_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1835 N_OUT9_Mn9@1835_d N_OUT8_Mn9@1835_g N_VSS_Mn9@1835_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1834 N_OUT9_Mn9@1834_d N_OUT8_Mn9@1834_g N_VSS_Mn9@1834_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1835 N_OUT9_Mp9@1835_d N_OUT8_Mp9@1835_g N_VDD_Mp9@1835_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1834 N_OUT9_Mp9@1834_d N_OUT8_Mp9@1834_g N_VDD_Mp9@1834_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1833 N_OUT9_Mn9@1833_d N_OUT8_Mn9@1833_g N_VSS_Mn9@1833_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1832 N_OUT9_Mn9@1832_d N_OUT8_Mn9@1832_g N_VSS_Mn9@1832_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1833 N_OUT9_Mp9@1833_d N_OUT8_Mp9@1833_g N_VDD_Mp9@1833_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1832 N_OUT9_Mp9@1832_d N_OUT8_Mp9@1832_g N_VDD_Mp9@1832_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1831 N_OUT9_Mn9@1831_d N_OUT8_Mn9@1831_g N_VSS_Mn9@1831_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1830 N_OUT9_Mn9@1830_d N_OUT8_Mn9@1830_g N_VSS_Mn9@1830_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1831 N_OUT9_Mp9@1831_d N_OUT8_Mp9@1831_g N_VDD_Mp9@1831_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1830 N_OUT9_Mp9@1830_d N_OUT8_Mp9@1830_g N_VDD_Mp9@1830_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1829 N_OUT9_Mn9@1829_d N_OUT8_Mn9@1829_g N_VSS_Mn9@1829_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1828 N_OUT9_Mn9@1828_d N_OUT8_Mn9@1828_g N_VSS_Mn9@1828_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1829 N_OUT9_Mp9@1829_d N_OUT8_Mp9@1829_g N_VDD_Mp9@1829_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1828 N_OUT9_Mp9@1828_d N_OUT8_Mp9@1828_g N_VDD_Mp9@1828_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1827 N_OUT9_Mn9@1827_d N_OUT8_Mn9@1827_g N_VSS_Mn9@1827_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1826 N_OUT9_Mn9@1826_d N_OUT8_Mn9@1826_g N_VSS_Mn9@1826_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1827 N_OUT9_Mp9@1827_d N_OUT8_Mp9@1827_g N_VDD_Mp9@1827_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1826 N_OUT9_Mp9@1826_d N_OUT8_Mp9@1826_g N_VDD_Mp9@1826_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1825 N_OUT9_Mn9@1825_d N_OUT8_Mn9@1825_g N_VSS_Mn9@1825_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1824 N_OUT9_Mn9@1824_d N_OUT8_Mn9@1824_g N_VSS_Mn9@1824_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1825 N_OUT9_Mp9@1825_d N_OUT8_Mp9@1825_g N_VDD_Mp9@1825_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1824 N_OUT9_Mp9@1824_d N_OUT8_Mp9@1824_g N_VDD_Mp9@1824_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1823 N_OUT9_Mn9@1823_d N_OUT8_Mn9@1823_g N_VSS_Mn9@1823_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1822 N_OUT9_Mn9@1822_d N_OUT8_Mn9@1822_g N_VSS_Mn9@1822_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1823 N_OUT9_Mp9@1823_d N_OUT8_Mp9@1823_g N_VDD_Mp9@1823_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1822 N_OUT9_Mp9@1822_d N_OUT8_Mp9@1822_g N_VDD_Mp9@1822_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1821 N_OUT9_Mn9@1821_d N_OUT8_Mn9@1821_g N_VSS_Mn9@1821_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1820 N_OUT9_Mn9@1820_d N_OUT8_Mn9@1820_g N_VSS_Mn9@1820_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1821 N_OUT9_Mp9@1821_d N_OUT8_Mp9@1821_g N_VDD_Mp9@1821_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1820 N_OUT9_Mp9@1820_d N_OUT8_Mp9@1820_g N_VDD_Mp9@1820_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1819 N_OUT9_Mn9@1819_d N_OUT8_Mn9@1819_g N_VSS_Mn9@1819_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1818 N_OUT9_Mn9@1818_d N_OUT8_Mn9@1818_g N_VSS_Mn9@1818_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1819 N_OUT9_Mp9@1819_d N_OUT8_Mp9@1819_g N_VDD_Mp9@1819_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1818 N_OUT9_Mp9@1818_d N_OUT8_Mp9@1818_g N_VDD_Mp9@1818_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1817 N_OUT9_Mn9@1817_d N_OUT8_Mn9@1817_g N_VSS_Mn9@1817_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1816 N_OUT9_Mn9@1816_d N_OUT8_Mn9@1816_g N_VSS_Mn9@1816_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1817 N_OUT9_Mp9@1817_d N_OUT8_Mp9@1817_g N_VDD_Mp9@1817_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1816 N_OUT9_Mp9@1816_d N_OUT8_Mp9@1816_g N_VDD_Mp9@1816_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1815 N_OUT9_Mn9@1815_d N_OUT8_Mn9@1815_g N_VSS_Mn9@1815_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1814 N_OUT9_Mn9@1814_d N_OUT8_Mn9@1814_g N_VSS_Mn9@1814_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1815 N_OUT9_Mp9@1815_d N_OUT8_Mp9@1815_g N_VDD_Mp9@1815_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1814 N_OUT9_Mp9@1814_d N_OUT8_Mp9@1814_g N_VDD_Mp9@1814_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1813 N_OUT9_Mn9@1813_d N_OUT8_Mn9@1813_g N_VSS_Mn9@1813_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1812 N_OUT9_Mn9@1812_d N_OUT8_Mn9@1812_g N_VSS_Mn9@1812_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1813 N_OUT9_Mp9@1813_d N_OUT8_Mp9@1813_g N_VDD_Mp9@1813_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1812 N_OUT9_Mp9@1812_d N_OUT8_Mp9@1812_g N_VDD_Mp9@1812_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1811 N_OUT9_Mn9@1811_d N_OUT8_Mn9@1811_g N_VSS_Mn9@1811_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1810 N_OUT9_Mn9@1810_d N_OUT8_Mn9@1810_g N_VSS_Mn9@1810_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1811 N_OUT9_Mp9@1811_d N_OUT8_Mp9@1811_g N_VDD_Mp9@1811_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1810 N_OUT9_Mp9@1810_d N_OUT8_Mp9@1810_g N_VDD_Mp9@1810_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1809 N_OUT9_Mn9@1809_d N_OUT8_Mn9@1809_g N_VSS_Mn9@1809_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1808 N_OUT9_Mn9@1808_d N_OUT8_Mn9@1808_g N_VSS_Mn9@1808_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1809 N_OUT9_Mp9@1809_d N_OUT8_Mp9@1809_g N_VDD_Mp9@1809_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1808 N_OUT9_Mp9@1808_d N_OUT8_Mp9@1808_g N_VDD_Mp9@1808_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1807 N_OUT9_Mn9@1807_d N_OUT8_Mn9@1807_g N_VSS_Mn9@1807_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1806 N_OUT9_Mn9@1806_d N_OUT8_Mn9@1806_g N_VSS_Mn9@1806_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1807 N_OUT9_Mp9@1807_d N_OUT8_Mp9@1807_g N_VDD_Mp9@1807_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1806 N_OUT9_Mp9@1806_d N_OUT8_Mp9@1806_g N_VDD_Mp9@1806_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1805 N_OUT9_Mn9@1805_d N_OUT8_Mn9@1805_g N_VSS_Mn9@1805_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1804 N_OUT9_Mn9@1804_d N_OUT8_Mn9@1804_g N_VSS_Mn9@1804_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1805 N_OUT9_Mp9@1805_d N_OUT8_Mp9@1805_g N_VDD_Mp9@1805_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1804 N_OUT9_Mp9@1804_d N_OUT8_Mp9@1804_g N_VDD_Mp9@1804_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1803 N_OUT9_Mn9@1803_d N_OUT8_Mn9@1803_g N_VSS_Mn9@1803_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1802 N_OUT9_Mn9@1802_d N_OUT8_Mn9@1802_g N_VSS_Mn9@1802_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1803 N_OUT9_Mp9@1803_d N_OUT8_Mp9@1803_g N_VDD_Mp9@1803_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1802 N_OUT9_Mp9@1802_d N_OUT8_Mp9@1802_g N_VDD_Mp9@1802_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1801 N_OUT9_Mn9@1801_d N_OUT8_Mn9@1801_g N_VSS_Mn9@1801_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1800 N_OUT9_Mn9@1800_d N_OUT8_Mn9@1800_g N_VSS_Mn9@1800_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1801 N_OUT9_Mp9@1801_d N_OUT8_Mp9@1801_g N_VDD_Mp9@1801_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1800 N_OUT9_Mp9@1800_d N_OUT8_Mp9@1800_g N_VDD_Mp9@1800_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1799 N_OUT9_Mn9@1799_d N_OUT8_Mn9@1799_g N_VSS_Mn9@1799_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1798 N_OUT9_Mn9@1798_d N_OUT8_Mn9@1798_g N_VSS_Mn9@1798_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1799 N_OUT9_Mp9@1799_d N_OUT8_Mp9@1799_g N_VDD_Mp9@1799_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1798 N_OUT9_Mp9@1798_d N_OUT8_Mp9@1798_g N_VDD_Mp9@1798_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1797 N_OUT9_Mn9@1797_d N_OUT8_Mn9@1797_g N_VSS_Mn9@1797_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1796 N_OUT9_Mn9@1796_d N_OUT8_Mn9@1796_g N_VSS_Mn9@1796_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1797 N_OUT9_Mp9@1797_d N_OUT8_Mp9@1797_g N_VDD_Mp9@1797_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1796 N_OUT9_Mp9@1796_d N_OUT8_Mp9@1796_g N_VDD_Mp9@1796_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1795 N_OUT9_Mn9@1795_d N_OUT8_Mn9@1795_g N_VSS_Mn9@1795_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1794 N_OUT9_Mn9@1794_d N_OUT8_Mn9@1794_g N_VSS_Mn9@1794_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1795 N_OUT9_Mp9@1795_d N_OUT8_Mp9@1795_g N_VDD_Mp9@1795_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1794 N_OUT9_Mp9@1794_d N_OUT8_Mp9@1794_g N_VDD_Mp9@1794_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1793 N_OUT9_Mn9@1793_d N_OUT8_Mn9@1793_g N_VSS_Mn9@1793_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1792 N_OUT9_Mn9@1792_d N_OUT8_Mn9@1792_g N_VSS_Mn9@1792_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1793 N_OUT9_Mp9@1793_d N_OUT8_Mp9@1793_g N_VDD_Mp9@1793_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1792 N_OUT9_Mp9@1792_d N_OUT8_Mp9@1792_g N_VDD_Mp9@1792_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1791 N_OUT9_Mn9@1791_d N_OUT8_Mn9@1791_g N_VSS_Mn9@1791_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1790 N_OUT9_Mn9@1790_d N_OUT8_Mn9@1790_g N_VSS_Mn9@1790_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1791 N_OUT9_Mp9@1791_d N_OUT8_Mp9@1791_g N_VDD_Mp9@1791_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1790 N_OUT9_Mp9@1790_d N_OUT8_Mp9@1790_g N_VDD_Mp9@1790_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1789 N_OUT9_Mn9@1789_d N_OUT8_Mn9@1789_g N_VSS_Mn9@1789_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1788 N_OUT9_Mn9@1788_d N_OUT8_Mn9@1788_g N_VSS_Mn9@1788_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1789 N_OUT9_Mp9@1789_d N_OUT8_Mp9@1789_g N_VDD_Mp9@1789_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1788 N_OUT9_Mp9@1788_d N_OUT8_Mp9@1788_g N_VDD_Mp9@1788_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1787 N_OUT9_Mn9@1787_d N_OUT8_Mn9@1787_g N_VSS_Mn9@1787_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1786 N_OUT9_Mn9@1786_d N_OUT8_Mn9@1786_g N_VSS_Mn9@1786_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1787 N_OUT9_Mp9@1787_d N_OUT8_Mp9@1787_g N_VDD_Mp9@1787_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1786 N_OUT9_Mp9@1786_d N_OUT8_Mp9@1786_g N_VDD_Mp9@1786_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1785 N_OUT9_Mn9@1785_d N_OUT8_Mn9@1785_g N_VSS_Mn9@1785_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1784 N_OUT9_Mn9@1784_d N_OUT8_Mn9@1784_g N_VSS_Mn9@1784_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1785 N_OUT9_Mp9@1785_d N_OUT8_Mp9@1785_g N_VDD_Mp9@1785_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1784 N_OUT9_Mp9@1784_d N_OUT8_Mp9@1784_g N_VDD_Mp9@1784_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1783 N_OUT9_Mn9@1783_d N_OUT8_Mn9@1783_g N_VSS_Mn9@1783_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1782 N_OUT9_Mn9@1782_d N_OUT8_Mn9@1782_g N_VSS_Mn9@1782_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1783 N_OUT9_Mp9@1783_d N_OUT8_Mp9@1783_g N_VDD_Mp9@1783_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1782 N_OUT9_Mp9@1782_d N_OUT8_Mp9@1782_g N_VDD_Mp9@1782_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1781 N_OUT9_Mn9@1781_d N_OUT8_Mn9@1781_g N_VSS_Mn9@1781_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1780 N_OUT9_Mn9@1780_d N_OUT8_Mn9@1780_g N_VSS_Mn9@1780_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1781 N_OUT9_Mp9@1781_d N_OUT8_Mp9@1781_g N_VDD_Mp9@1781_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1780 N_OUT9_Mp9@1780_d N_OUT8_Mp9@1780_g N_VDD_Mp9@1780_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1779 N_OUT9_Mn9@1779_d N_OUT8_Mn9@1779_g N_VSS_Mn9@1779_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1778 N_OUT9_Mn9@1778_d N_OUT8_Mn9@1778_g N_VSS_Mn9@1778_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1779 N_OUT9_Mp9@1779_d N_OUT8_Mp9@1779_g N_VDD_Mp9@1779_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1778 N_OUT9_Mp9@1778_d N_OUT8_Mp9@1778_g N_VDD_Mp9@1778_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1777 N_OUT9_Mn9@1777_d N_OUT8_Mn9@1777_g N_VSS_Mn9@1777_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1776 N_OUT9_Mn9@1776_d N_OUT8_Mn9@1776_g N_VSS_Mn9@1776_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1777 N_OUT9_Mp9@1777_d N_OUT8_Mp9@1777_g N_VDD_Mp9@1777_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1776 N_OUT9_Mp9@1776_d N_OUT8_Mp9@1776_g N_VDD_Mp9@1776_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1775 N_OUT9_Mn9@1775_d N_OUT8_Mn9@1775_g N_VSS_Mn9@1775_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1774 N_OUT9_Mn9@1774_d N_OUT8_Mn9@1774_g N_VSS_Mn9@1774_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1775 N_OUT9_Mp9@1775_d N_OUT8_Mp9@1775_g N_VDD_Mp9@1775_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1774 N_OUT9_Mp9@1774_d N_OUT8_Mp9@1774_g N_VDD_Mp9@1774_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1773 N_OUT9_Mn9@1773_d N_OUT8_Mn9@1773_g N_VSS_Mn9@1773_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1772 N_OUT9_Mn9@1772_d N_OUT8_Mn9@1772_g N_VSS_Mn9@1772_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1773 N_OUT9_Mp9@1773_d N_OUT8_Mp9@1773_g N_VDD_Mp9@1773_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1772 N_OUT9_Mp9@1772_d N_OUT8_Mp9@1772_g N_VDD_Mp9@1772_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1771 N_OUT9_Mn9@1771_d N_OUT8_Mn9@1771_g N_VSS_Mn9@1771_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1770 N_OUT9_Mn9@1770_d N_OUT8_Mn9@1770_g N_VSS_Mn9@1770_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1771 N_OUT9_Mp9@1771_d N_OUT8_Mp9@1771_g N_VDD_Mp9@1771_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1770 N_OUT9_Mp9@1770_d N_OUT8_Mp9@1770_g N_VDD_Mp9@1770_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1769 N_OUT9_Mn9@1769_d N_OUT8_Mn9@1769_g N_VSS_Mn9@1769_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1768 N_OUT9_Mn9@1768_d N_OUT8_Mn9@1768_g N_VSS_Mn9@1768_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1769 N_OUT9_Mp9@1769_d N_OUT8_Mp9@1769_g N_VDD_Mp9@1769_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1768 N_OUT9_Mp9@1768_d N_OUT8_Mp9@1768_g N_VDD_Mp9@1768_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1767 N_OUT9_Mn9@1767_d N_OUT8_Mn9@1767_g N_VSS_Mn9@1767_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1766 N_OUT9_Mn9@1766_d N_OUT8_Mn9@1766_g N_VSS_Mn9@1766_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1767 N_OUT9_Mp9@1767_d N_OUT8_Mp9@1767_g N_VDD_Mp9@1767_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1766 N_OUT9_Mp9@1766_d N_OUT8_Mp9@1766_g N_VDD_Mp9@1766_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1765 N_OUT9_Mn9@1765_d N_OUT8_Mn9@1765_g N_VSS_Mn9@1765_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1764 N_OUT9_Mn9@1764_d N_OUT8_Mn9@1764_g N_VSS_Mn9@1764_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1765 N_OUT9_Mp9@1765_d N_OUT8_Mp9@1765_g N_VDD_Mp9@1765_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1764 N_OUT9_Mp9@1764_d N_OUT8_Mp9@1764_g N_VDD_Mp9@1764_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1763 N_OUT9_Mn9@1763_d N_OUT8_Mn9@1763_g N_VSS_Mn9@1763_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1762 N_OUT9_Mn9@1762_d N_OUT8_Mn9@1762_g N_VSS_Mn9@1762_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1763 N_OUT9_Mp9@1763_d N_OUT8_Mp9@1763_g N_VDD_Mp9@1763_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1762 N_OUT9_Mp9@1762_d N_OUT8_Mp9@1762_g N_VDD_Mp9@1762_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1761 N_OUT9_Mn9@1761_d N_OUT8_Mn9@1761_g N_VSS_Mn9@1761_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1760 N_OUT9_Mn9@1760_d N_OUT8_Mn9@1760_g N_VSS_Mn9@1760_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1761 N_OUT9_Mp9@1761_d N_OUT8_Mp9@1761_g N_VDD_Mp9@1761_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1760 N_OUT9_Mp9@1760_d N_OUT8_Mp9@1760_g N_VDD_Mp9@1760_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1759 N_OUT9_Mn9@1759_d N_OUT8_Mn9@1759_g N_VSS_Mn9@1759_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1758 N_OUT9_Mn9@1758_d N_OUT8_Mn9@1758_g N_VSS_Mn9@1758_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1759 N_OUT9_Mp9@1759_d N_OUT8_Mp9@1759_g N_VDD_Mp9@1759_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1758 N_OUT9_Mp9@1758_d N_OUT8_Mp9@1758_g N_VDD_Mp9@1758_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1757 N_OUT9_Mn9@1757_d N_OUT8_Mn9@1757_g N_VSS_Mn9@1757_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1756 N_OUT9_Mn9@1756_d N_OUT8_Mn9@1756_g N_VSS_Mn9@1756_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1757 N_OUT9_Mp9@1757_d N_OUT8_Mp9@1757_g N_VDD_Mp9@1757_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1756 N_OUT9_Mp9@1756_d N_OUT8_Mp9@1756_g N_VDD_Mp9@1756_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1755 N_OUT9_Mn9@1755_d N_OUT8_Mn9@1755_g N_VSS_Mn9@1755_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1754 N_OUT9_Mn9@1754_d N_OUT8_Mn9@1754_g N_VSS_Mn9@1754_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1755 N_OUT9_Mp9@1755_d N_OUT8_Mp9@1755_g N_VDD_Mp9@1755_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1754 N_OUT9_Mp9@1754_d N_OUT8_Mp9@1754_g N_VDD_Mp9@1754_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1753 N_OUT9_Mn9@1753_d N_OUT8_Mn9@1753_g N_VSS_Mn9@1753_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1752 N_OUT9_Mn9@1752_d N_OUT8_Mn9@1752_g N_VSS_Mn9@1752_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1753 N_OUT9_Mp9@1753_d N_OUT8_Mp9@1753_g N_VDD_Mp9@1753_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1752 N_OUT9_Mp9@1752_d N_OUT8_Mp9@1752_g N_VDD_Mp9@1752_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1751 N_OUT9_Mn9@1751_d N_OUT8_Mn9@1751_g N_VSS_Mn9@1751_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1750 N_OUT9_Mn9@1750_d N_OUT8_Mn9@1750_g N_VSS_Mn9@1750_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1751 N_OUT9_Mp9@1751_d N_OUT8_Mp9@1751_g N_VDD_Mp9@1751_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1750 N_OUT9_Mp9@1750_d N_OUT8_Mp9@1750_g N_VDD_Mp9@1750_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1749 N_OUT9_Mn9@1749_d N_OUT8_Mn9@1749_g N_VSS_Mn9@1749_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1748 N_OUT9_Mn9@1748_d N_OUT8_Mn9@1748_g N_VSS_Mn9@1748_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1749 N_OUT9_Mp9@1749_d N_OUT8_Mp9@1749_g N_VDD_Mp9@1749_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1748 N_OUT9_Mp9@1748_d N_OUT8_Mp9@1748_g N_VDD_Mp9@1748_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1747 N_OUT9_Mn9@1747_d N_OUT8_Mn9@1747_g N_VSS_Mn9@1747_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1746 N_OUT9_Mn9@1746_d N_OUT8_Mn9@1746_g N_VSS_Mn9@1746_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1747 N_OUT9_Mp9@1747_d N_OUT8_Mp9@1747_g N_VDD_Mp9@1747_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1746 N_OUT9_Mp9@1746_d N_OUT8_Mp9@1746_g N_VDD_Mp9@1746_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1745 N_OUT9_Mn9@1745_d N_OUT8_Mn9@1745_g N_VSS_Mn9@1745_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1744 N_OUT9_Mn9@1744_d N_OUT8_Mn9@1744_g N_VSS_Mn9@1744_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1745 N_OUT9_Mp9@1745_d N_OUT8_Mp9@1745_g N_VDD_Mp9@1745_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1744 N_OUT9_Mp9@1744_d N_OUT8_Mp9@1744_g N_VDD_Mp9@1744_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1743 N_OUT9_Mn9@1743_d N_OUT8_Mn9@1743_g N_VSS_Mn9@1743_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1742 N_OUT9_Mn9@1742_d N_OUT8_Mn9@1742_g N_VSS_Mn9@1742_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1743 N_OUT9_Mp9@1743_d N_OUT8_Mp9@1743_g N_VDD_Mp9@1743_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1742 N_OUT9_Mp9@1742_d N_OUT8_Mp9@1742_g N_VDD_Mp9@1742_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1741 N_OUT9_Mn9@1741_d N_OUT8_Mn9@1741_g N_VSS_Mn9@1741_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1740 N_OUT9_Mn9@1740_d N_OUT8_Mn9@1740_g N_VSS_Mn9@1740_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1741 N_OUT9_Mp9@1741_d N_OUT8_Mp9@1741_g N_VDD_Mp9@1741_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1740 N_OUT9_Mp9@1740_d N_OUT8_Mp9@1740_g N_VDD_Mp9@1740_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1739 N_OUT9_Mn9@1739_d N_OUT8_Mn9@1739_g N_VSS_Mn9@1739_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1738 N_OUT9_Mn9@1738_d N_OUT8_Mn9@1738_g N_VSS_Mn9@1738_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1739 N_OUT9_Mp9@1739_d N_OUT8_Mp9@1739_g N_VDD_Mp9@1739_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1738 N_OUT9_Mp9@1738_d N_OUT8_Mp9@1738_g N_VDD_Mp9@1738_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1737 N_OUT9_Mn9@1737_d N_OUT8_Mn9@1737_g N_VSS_Mn9@1737_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1736 N_OUT9_Mn9@1736_d N_OUT8_Mn9@1736_g N_VSS_Mn9@1736_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1737 N_OUT9_Mp9@1737_d N_OUT8_Mp9@1737_g N_VDD_Mp9@1737_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1736 N_OUT9_Mp9@1736_d N_OUT8_Mp9@1736_g N_VDD_Mp9@1736_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1735 N_OUT9_Mn9@1735_d N_OUT8_Mn9@1735_g N_VSS_Mn9@1735_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1734 N_OUT9_Mn9@1734_d N_OUT8_Mn9@1734_g N_VSS_Mn9@1734_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1735 N_OUT9_Mp9@1735_d N_OUT8_Mp9@1735_g N_VDD_Mp9@1735_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1734 N_OUT9_Mp9@1734_d N_OUT8_Mp9@1734_g N_VDD_Mp9@1734_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1733 N_OUT9_Mn9@1733_d N_OUT8_Mn9@1733_g N_VSS_Mn9@1733_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1732 N_OUT9_Mn9@1732_d N_OUT8_Mn9@1732_g N_VSS_Mn9@1732_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1733 N_OUT9_Mp9@1733_d N_OUT8_Mp9@1733_g N_VDD_Mp9@1733_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1732 N_OUT9_Mp9@1732_d N_OUT8_Mp9@1732_g N_VDD_Mp9@1732_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1731 N_OUT9_Mn9@1731_d N_OUT8_Mn9@1731_g N_VSS_Mn9@1731_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1730 N_OUT9_Mn9@1730_d N_OUT8_Mn9@1730_g N_VSS_Mn9@1730_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1731 N_OUT9_Mp9@1731_d N_OUT8_Mp9@1731_g N_VDD_Mp9@1731_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1730 N_OUT9_Mp9@1730_d N_OUT8_Mp9@1730_g N_VDD_Mp9@1730_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1729 N_OUT9_Mn9@1729_d N_OUT8_Mn9@1729_g N_VSS_Mn9@1729_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1728 N_OUT9_Mn9@1728_d N_OUT8_Mn9@1728_g N_VSS_Mn9@1728_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1729 N_OUT9_Mp9@1729_d N_OUT8_Mp9@1729_g N_VDD_Mp9@1729_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1728 N_OUT9_Mp9@1728_d N_OUT8_Mp9@1728_g N_VDD_Mp9@1728_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1727 N_OUT9_Mn9@1727_d N_OUT8_Mn9@1727_g N_VSS_Mn9@1727_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1726 N_OUT9_Mn9@1726_d N_OUT8_Mn9@1726_g N_VSS_Mn9@1726_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1727 N_OUT9_Mp9@1727_d N_OUT8_Mp9@1727_g N_VDD_Mp9@1727_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1726 N_OUT9_Mp9@1726_d N_OUT8_Mp9@1726_g N_VDD_Mp9@1726_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1725 N_OUT9_Mn9@1725_d N_OUT8_Mn9@1725_g N_VSS_Mn9@1725_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1724 N_OUT9_Mn9@1724_d N_OUT8_Mn9@1724_g N_VSS_Mn9@1724_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1725 N_OUT9_Mp9@1725_d N_OUT8_Mp9@1725_g N_VDD_Mp9@1725_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1724 N_OUT9_Mp9@1724_d N_OUT8_Mp9@1724_g N_VDD_Mp9@1724_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1723 N_OUT9_Mn9@1723_d N_OUT8_Mn9@1723_g N_VSS_Mn9@1723_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1722 N_OUT9_Mn9@1722_d N_OUT8_Mn9@1722_g N_VSS_Mn9@1722_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1723 N_OUT9_Mp9@1723_d N_OUT8_Mp9@1723_g N_VDD_Mp9@1723_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1722 N_OUT9_Mp9@1722_d N_OUT8_Mp9@1722_g N_VDD_Mp9@1722_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1721 N_OUT9_Mn9@1721_d N_OUT8_Mn9@1721_g N_VSS_Mn9@1721_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1720 N_OUT9_Mn9@1720_d N_OUT8_Mn9@1720_g N_VSS_Mn9@1720_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1721 N_OUT9_Mp9@1721_d N_OUT8_Mp9@1721_g N_VDD_Mp9@1721_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1720 N_OUT9_Mp9@1720_d N_OUT8_Mp9@1720_g N_VDD_Mp9@1720_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1719 N_OUT9_Mn9@1719_d N_OUT8_Mn9@1719_g N_VSS_Mn9@1719_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1718 N_OUT9_Mn9@1718_d N_OUT8_Mn9@1718_g N_VSS_Mn9@1718_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1719 N_OUT9_Mp9@1719_d N_OUT8_Mp9@1719_g N_VDD_Mp9@1719_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1718 N_OUT9_Mp9@1718_d N_OUT8_Mp9@1718_g N_VDD_Mp9@1718_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1717 N_OUT9_Mn9@1717_d N_OUT8_Mn9@1717_g N_VSS_Mn9@1717_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1716 N_OUT9_Mn9@1716_d N_OUT8_Mn9@1716_g N_VSS_Mn9@1716_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1717 N_OUT9_Mp9@1717_d N_OUT8_Mp9@1717_g N_VDD_Mp9@1717_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1716 N_OUT9_Mp9@1716_d N_OUT8_Mp9@1716_g N_VDD_Mp9@1716_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1715 N_OUT9_Mn9@1715_d N_OUT8_Mn9@1715_g N_VSS_Mn9@1715_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1714 N_OUT9_Mn9@1714_d N_OUT8_Mn9@1714_g N_VSS_Mn9@1714_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1715 N_OUT9_Mp9@1715_d N_OUT8_Mp9@1715_g N_VDD_Mp9@1715_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1714 N_OUT9_Mp9@1714_d N_OUT8_Mp9@1714_g N_VDD_Mp9@1714_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1713 N_OUT9_Mn9@1713_d N_OUT8_Mn9@1713_g N_VSS_Mn9@1713_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1712 N_OUT9_Mn9@1712_d N_OUT8_Mn9@1712_g N_VSS_Mn9@1712_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1713 N_OUT9_Mp9@1713_d N_OUT8_Mp9@1713_g N_VDD_Mp9@1713_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1712 N_OUT9_Mp9@1712_d N_OUT8_Mp9@1712_g N_VDD_Mp9@1712_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1711 N_OUT9_Mn9@1711_d N_OUT8_Mn9@1711_g N_VSS_Mn9@1711_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1710 N_OUT9_Mn9@1710_d N_OUT8_Mn9@1710_g N_VSS_Mn9@1710_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1711 N_OUT9_Mp9@1711_d N_OUT8_Mp9@1711_g N_VDD_Mp9@1711_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1710 N_OUT9_Mp9@1710_d N_OUT8_Mp9@1710_g N_VDD_Mp9@1710_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1709 N_OUT9_Mn9@1709_d N_OUT8_Mn9@1709_g N_VSS_Mn9@1709_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1708 N_OUT9_Mn9@1708_d N_OUT8_Mn9@1708_g N_VSS_Mn9@1708_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1709 N_OUT9_Mp9@1709_d N_OUT8_Mp9@1709_g N_VDD_Mp9@1709_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1708 N_OUT9_Mp9@1708_d N_OUT8_Mp9@1708_g N_VDD_Mp9@1708_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1707 N_OUT9_Mn9@1707_d N_OUT8_Mn9@1707_g N_VSS_Mn9@1707_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1706 N_OUT9_Mn9@1706_d N_OUT8_Mn9@1706_g N_VSS_Mn9@1706_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1707 N_OUT9_Mp9@1707_d N_OUT8_Mp9@1707_g N_VDD_Mp9@1707_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1706 N_OUT9_Mp9@1706_d N_OUT8_Mp9@1706_g N_VDD_Mp9@1706_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1705 N_OUT9_Mn9@1705_d N_OUT8_Mn9@1705_g N_VSS_Mn9@1705_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1704 N_OUT9_Mn9@1704_d N_OUT8_Mn9@1704_g N_VSS_Mn9@1704_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1705 N_OUT9_Mp9@1705_d N_OUT8_Mp9@1705_g N_VDD_Mp9@1705_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1704 N_OUT9_Mp9@1704_d N_OUT8_Mp9@1704_g N_VDD_Mp9@1704_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1703 N_OUT9_Mn9@1703_d N_OUT8_Mn9@1703_g N_VSS_Mn9@1703_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1702 N_OUT9_Mn9@1702_d N_OUT8_Mn9@1702_g N_VSS_Mn9@1702_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1703 N_OUT9_Mp9@1703_d N_OUT8_Mp9@1703_g N_VDD_Mp9@1703_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1702 N_OUT9_Mp9@1702_d N_OUT8_Mp9@1702_g N_VDD_Mp9@1702_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1701 N_OUT9_Mn9@1701_d N_OUT8_Mn9@1701_g N_VSS_Mn9@1701_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1700 N_OUT9_Mn9@1700_d N_OUT8_Mn9@1700_g N_VSS_Mn9@1700_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1701 N_OUT9_Mp9@1701_d N_OUT8_Mp9@1701_g N_VDD_Mp9@1701_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1700 N_OUT9_Mp9@1700_d N_OUT8_Mp9@1700_g N_VDD_Mp9@1700_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1699 N_OUT9_Mn9@1699_d N_OUT8_Mn9@1699_g N_VSS_Mn9@1699_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1698 N_OUT9_Mn9@1698_d N_OUT8_Mn9@1698_g N_VSS_Mn9@1698_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1699 N_OUT9_Mp9@1699_d N_OUT8_Mp9@1699_g N_VDD_Mp9@1699_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1698 N_OUT9_Mp9@1698_d N_OUT8_Mp9@1698_g N_VDD_Mp9@1698_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1697 N_OUT9_Mn9@1697_d N_OUT8_Mn9@1697_g N_VSS_Mn9@1697_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1696 N_OUT9_Mn9@1696_d N_OUT8_Mn9@1696_g N_VSS_Mn9@1696_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1697 N_OUT9_Mp9@1697_d N_OUT8_Mp9@1697_g N_VDD_Mp9@1697_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1696 N_OUT9_Mp9@1696_d N_OUT8_Mp9@1696_g N_VDD_Mp9@1696_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1695 N_OUT9_Mn9@1695_d N_OUT8_Mn9@1695_g N_VSS_Mn9@1695_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1694 N_OUT9_Mn9@1694_d N_OUT8_Mn9@1694_g N_VSS_Mn9@1694_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1695 N_OUT9_Mp9@1695_d N_OUT8_Mp9@1695_g N_VDD_Mp9@1695_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1694 N_OUT9_Mp9@1694_d N_OUT8_Mp9@1694_g N_VDD_Mp9@1694_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1693 N_OUT9_Mn9@1693_d N_OUT8_Mn9@1693_g N_VSS_Mn9@1693_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1692 N_OUT9_Mn9@1692_d N_OUT8_Mn9@1692_g N_VSS_Mn9@1692_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1693 N_OUT9_Mp9@1693_d N_OUT8_Mp9@1693_g N_VDD_Mp9@1693_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1692 N_OUT9_Mp9@1692_d N_OUT8_Mp9@1692_g N_VDD_Mp9@1692_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1691 N_OUT9_Mn9@1691_d N_OUT8_Mn9@1691_g N_VSS_Mn9@1691_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1690 N_OUT9_Mn9@1690_d N_OUT8_Mn9@1690_g N_VSS_Mn9@1690_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1691 N_OUT9_Mp9@1691_d N_OUT8_Mp9@1691_g N_VDD_Mp9@1691_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1690 N_OUT9_Mp9@1690_d N_OUT8_Mp9@1690_g N_VDD_Mp9@1690_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1689 N_OUT9_Mn9@1689_d N_OUT8_Mn9@1689_g N_VSS_Mn9@1689_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1688 N_OUT9_Mn9@1688_d N_OUT8_Mn9@1688_g N_VSS_Mn9@1688_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1689 N_OUT9_Mp9@1689_d N_OUT8_Mp9@1689_g N_VDD_Mp9@1689_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1688 N_OUT9_Mp9@1688_d N_OUT8_Mp9@1688_g N_VDD_Mp9@1688_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1687 N_OUT9_Mn9@1687_d N_OUT8_Mn9@1687_g N_VSS_Mn9@1687_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1686 N_OUT9_Mn9@1686_d N_OUT8_Mn9@1686_g N_VSS_Mn9@1686_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1687 N_OUT9_Mp9@1687_d N_OUT8_Mp9@1687_g N_VDD_Mp9@1687_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1686 N_OUT9_Mp9@1686_d N_OUT8_Mp9@1686_g N_VDD_Mp9@1686_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1685 N_OUT9_Mn9@1685_d N_OUT8_Mn9@1685_g N_VSS_Mn9@1685_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1684 N_OUT9_Mn9@1684_d N_OUT8_Mn9@1684_g N_VSS_Mn9@1684_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1685 N_OUT9_Mp9@1685_d N_OUT8_Mp9@1685_g N_VDD_Mp9@1685_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1684 N_OUT9_Mp9@1684_d N_OUT8_Mp9@1684_g N_VDD_Mp9@1684_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1683 N_OUT9_Mn9@1683_d N_OUT8_Mn9@1683_g N_VSS_Mn9@1683_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1682 N_OUT9_Mn9@1682_d N_OUT8_Mn9@1682_g N_VSS_Mn9@1682_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1683 N_OUT9_Mp9@1683_d N_OUT8_Mp9@1683_g N_VDD_Mp9@1683_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1682 N_OUT9_Mp9@1682_d N_OUT8_Mp9@1682_g N_VDD_Mp9@1682_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1681 N_OUT9_Mn9@1681_d N_OUT8_Mn9@1681_g N_VSS_Mn9@1681_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1680 N_OUT9_Mn9@1680_d N_OUT8_Mn9@1680_g N_VSS_Mn9@1680_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1681 N_OUT9_Mp9@1681_d N_OUT8_Mp9@1681_g N_VDD_Mp9@1681_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1680 N_OUT9_Mp9@1680_d N_OUT8_Mp9@1680_g N_VDD_Mp9@1680_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1679 N_OUT9_Mn9@1679_d N_OUT8_Mn9@1679_g N_VSS_Mn9@1679_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1678 N_OUT9_Mn9@1678_d N_OUT8_Mn9@1678_g N_VSS_Mn9@1678_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1679 N_OUT9_Mp9@1679_d N_OUT8_Mp9@1679_g N_VDD_Mp9@1679_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1678 N_OUT9_Mp9@1678_d N_OUT8_Mp9@1678_g N_VDD_Mp9@1678_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1677 N_OUT9_Mn9@1677_d N_OUT8_Mn9@1677_g N_VSS_Mn9@1677_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1676 N_OUT9_Mn9@1676_d N_OUT8_Mn9@1676_g N_VSS_Mn9@1676_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1677 N_OUT9_Mp9@1677_d N_OUT8_Mp9@1677_g N_VDD_Mp9@1677_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1676 N_OUT9_Mp9@1676_d N_OUT8_Mp9@1676_g N_VDD_Mp9@1676_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1675 N_OUT9_Mn9@1675_d N_OUT8_Mn9@1675_g N_VSS_Mn9@1675_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1674 N_OUT9_Mn9@1674_d N_OUT8_Mn9@1674_g N_VSS_Mn9@1674_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1675 N_OUT9_Mp9@1675_d N_OUT8_Mp9@1675_g N_VDD_Mp9@1675_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1674 N_OUT9_Mp9@1674_d N_OUT8_Mp9@1674_g N_VDD_Mp9@1674_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1673 N_OUT9_Mn9@1673_d N_OUT8_Mn9@1673_g N_VSS_Mn9@1673_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1672 N_OUT9_Mn9@1672_d N_OUT8_Mn9@1672_g N_VSS_Mn9@1672_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1673 N_OUT9_Mp9@1673_d N_OUT8_Mp9@1673_g N_VDD_Mp9@1673_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1672 N_OUT9_Mp9@1672_d N_OUT8_Mp9@1672_g N_VDD_Mp9@1672_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1671 N_OUT9_Mn9@1671_d N_OUT8_Mn9@1671_g N_VSS_Mn9@1671_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1670 N_OUT9_Mn9@1670_d N_OUT8_Mn9@1670_g N_VSS_Mn9@1670_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1671 N_OUT9_Mp9@1671_d N_OUT8_Mp9@1671_g N_VDD_Mp9@1671_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1670 N_OUT9_Mp9@1670_d N_OUT8_Mp9@1670_g N_VDD_Mp9@1670_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1669 N_OUT9_Mn9@1669_d N_OUT8_Mn9@1669_g N_VSS_Mn9@1669_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1668 N_OUT9_Mn9@1668_d N_OUT8_Mn9@1668_g N_VSS_Mn9@1668_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1669 N_OUT9_Mp9@1669_d N_OUT8_Mp9@1669_g N_VDD_Mp9@1669_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1668 N_OUT9_Mp9@1668_d N_OUT8_Mp9@1668_g N_VDD_Mp9@1668_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1667 N_OUT9_Mn9@1667_d N_OUT8_Mn9@1667_g N_VSS_Mn9@1667_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1666 N_OUT9_Mn9@1666_d N_OUT8_Mn9@1666_g N_VSS_Mn9@1666_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1667 N_OUT9_Mp9@1667_d N_OUT8_Mp9@1667_g N_VDD_Mp9@1667_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1666 N_OUT9_Mp9@1666_d N_OUT8_Mp9@1666_g N_VDD_Mp9@1666_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1665 N_OUT9_Mn9@1665_d N_OUT8_Mn9@1665_g N_VSS_Mn9@1665_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1664 N_OUT9_Mn9@1664_d N_OUT8_Mn9@1664_g N_VSS_Mn9@1664_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1665 N_OUT9_Mp9@1665_d N_OUT8_Mp9@1665_g N_VDD_Mp9@1665_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1664 N_OUT9_Mp9@1664_d N_OUT8_Mp9@1664_g N_VDD_Mp9@1664_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1663 N_OUT9_Mn9@1663_d N_OUT8_Mn9@1663_g N_VSS_Mn9@1663_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1662 N_OUT9_Mn9@1662_d N_OUT8_Mn9@1662_g N_VSS_Mn9@1662_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1663 N_OUT9_Mp9@1663_d N_OUT8_Mp9@1663_g N_VDD_Mp9@1663_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1662 N_OUT9_Mp9@1662_d N_OUT8_Mp9@1662_g N_VDD_Mp9@1662_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1661 N_OUT9_Mn9@1661_d N_OUT8_Mn9@1661_g N_VSS_Mn9@1661_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1660 N_OUT9_Mn9@1660_d N_OUT8_Mn9@1660_g N_VSS_Mn9@1660_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1661 N_OUT9_Mp9@1661_d N_OUT8_Mp9@1661_g N_VDD_Mp9@1661_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1660 N_OUT9_Mp9@1660_d N_OUT8_Mp9@1660_g N_VDD_Mp9@1660_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1659 N_OUT9_Mn9@1659_d N_OUT8_Mn9@1659_g N_VSS_Mn9@1659_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1658 N_OUT9_Mn9@1658_d N_OUT8_Mn9@1658_g N_VSS_Mn9@1658_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1659 N_OUT9_Mp9@1659_d N_OUT8_Mp9@1659_g N_VDD_Mp9@1659_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1658 N_OUT9_Mp9@1658_d N_OUT8_Mp9@1658_g N_VDD_Mp9@1658_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1657 N_OUT9_Mn9@1657_d N_OUT8_Mn9@1657_g N_VSS_Mn9@1657_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1656 N_OUT9_Mn9@1656_d N_OUT8_Mn9@1656_g N_VSS_Mn9@1656_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1657 N_OUT9_Mp9@1657_d N_OUT8_Mp9@1657_g N_VDD_Mp9@1657_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1656 N_OUT9_Mp9@1656_d N_OUT8_Mp9@1656_g N_VDD_Mp9@1656_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1655 N_OUT9_Mn9@1655_d N_OUT8_Mn9@1655_g N_VSS_Mn9@1655_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1654 N_OUT9_Mn9@1654_d N_OUT8_Mn9@1654_g N_VSS_Mn9@1654_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1655 N_OUT9_Mp9@1655_d N_OUT8_Mp9@1655_g N_VDD_Mp9@1655_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1654 N_OUT9_Mp9@1654_d N_OUT8_Mp9@1654_g N_VDD_Mp9@1654_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1653 N_OUT9_Mn9@1653_d N_OUT8_Mn9@1653_g N_VSS_Mn9@1653_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1652 N_OUT9_Mn9@1652_d N_OUT8_Mn9@1652_g N_VSS_Mn9@1652_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1653 N_OUT9_Mp9@1653_d N_OUT8_Mp9@1653_g N_VDD_Mp9@1653_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1652 N_OUT9_Mp9@1652_d N_OUT8_Mp9@1652_g N_VDD_Mp9@1652_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1651 N_OUT9_Mn9@1651_d N_OUT8_Mn9@1651_g N_VSS_Mn9@1651_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1650 N_OUT9_Mn9@1650_d N_OUT8_Mn9@1650_g N_VSS_Mn9@1650_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1651 N_OUT9_Mp9@1651_d N_OUT8_Mp9@1651_g N_VDD_Mp9@1651_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1650 N_OUT9_Mp9@1650_d N_OUT8_Mp9@1650_g N_VDD_Mp9@1650_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1649 N_OUT9_Mn9@1649_d N_OUT8_Mn9@1649_g N_VSS_Mn9@1649_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1648 N_OUT9_Mn9@1648_d N_OUT8_Mn9@1648_g N_VSS_Mn9@1648_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1649 N_OUT9_Mp9@1649_d N_OUT8_Mp9@1649_g N_VDD_Mp9@1649_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1648 N_OUT9_Mp9@1648_d N_OUT8_Mp9@1648_g N_VDD_Mp9@1648_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1647 N_OUT9_Mn9@1647_d N_OUT8_Mn9@1647_g N_VSS_Mn9@1647_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1646 N_OUT9_Mn9@1646_d N_OUT8_Mn9@1646_g N_VSS_Mn9@1646_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1647 N_OUT9_Mp9@1647_d N_OUT8_Mp9@1647_g N_VDD_Mp9@1647_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1646 N_OUT9_Mp9@1646_d N_OUT8_Mp9@1646_g N_VDD_Mp9@1646_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1645 N_OUT9_Mn9@1645_d N_OUT8_Mn9@1645_g N_VSS_Mn9@1645_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1644 N_OUT9_Mn9@1644_d N_OUT8_Mn9@1644_g N_VSS_Mn9@1644_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1645 N_OUT9_Mp9@1645_d N_OUT8_Mp9@1645_g N_VDD_Mp9@1645_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1644 N_OUT9_Mp9@1644_d N_OUT8_Mp9@1644_g N_VDD_Mp9@1644_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1643 N_OUT9_Mn9@1643_d N_OUT8_Mn9@1643_g N_VSS_Mn9@1643_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1642 N_OUT9_Mn9@1642_d N_OUT8_Mn9@1642_g N_VSS_Mn9@1642_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1643 N_OUT9_Mp9@1643_d N_OUT8_Mp9@1643_g N_VDD_Mp9@1643_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1642 N_OUT9_Mp9@1642_d N_OUT8_Mp9@1642_g N_VDD_Mp9@1642_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1641 N_OUT9_Mn9@1641_d N_OUT8_Mn9@1641_g N_VSS_Mn9@1641_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1640 N_OUT9_Mn9@1640_d N_OUT8_Mn9@1640_g N_VSS_Mn9@1640_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1641 N_OUT9_Mp9@1641_d N_OUT8_Mp9@1641_g N_VDD_Mp9@1641_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1640 N_OUT9_Mp9@1640_d N_OUT8_Mp9@1640_g N_VDD_Mp9@1640_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1639 N_OUT9_Mn9@1639_d N_OUT8_Mn9@1639_g N_VSS_Mn9@1639_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1638 N_OUT9_Mn9@1638_d N_OUT8_Mn9@1638_g N_VSS_Mn9@1638_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1639 N_OUT9_Mp9@1639_d N_OUT8_Mp9@1639_g N_VDD_Mp9@1639_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1638 N_OUT9_Mp9@1638_d N_OUT8_Mp9@1638_g N_VDD_Mp9@1638_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1637 N_OUT9_Mn9@1637_d N_OUT8_Mn9@1637_g N_VSS_Mn9@1637_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1636 N_OUT9_Mn9@1636_d N_OUT8_Mn9@1636_g N_VSS_Mn9@1636_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1637 N_OUT9_Mp9@1637_d N_OUT8_Mp9@1637_g N_VDD_Mp9@1637_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1636 N_OUT9_Mp9@1636_d N_OUT8_Mp9@1636_g N_VDD_Mp9@1636_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1635 N_OUT9_Mn9@1635_d N_OUT8_Mn9@1635_g N_VSS_Mn9@1635_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1634 N_OUT9_Mn9@1634_d N_OUT8_Mn9@1634_g N_VSS_Mn9@1634_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1635 N_OUT9_Mp9@1635_d N_OUT8_Mp9@1635_g N_VDD_Mp9@1635_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1634 N_OUT9_Mp9@1634_d N_OUT8_Mp9@1634_g N_VDD_Mp9@1634_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1633 N_OUT9_Mn9@1633_d N_OUT8_Mn9@1633_g N_VSS_Mn9@1633_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1632 N_OUT9_Mn9@1632_d N_OUT8_Mn9@1632_g N_VSS_Mn9@1632_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1633 N_OUT9_Mp9@1633_d N_OUT8_Mp9@1633_g N_VDD_Mp9@1633_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1632 N_OUT9_Mp9@1632_d N_OUT8_Mp9@1632_g N_VDD_Mp9@1632_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1631 N_OUT9_Mn9@1631_d N_OUT8_Mn9@1631_g N_VSS_Mn9@1631_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1630 N_OUT9_Mn9@1630_d N_OUT8_Mn9@1630_g N_VSS_Mn9@1630_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1631 N_OUT9_Mp9@1631_d N_OUT8_Mp9@1631_g N_VDD_Mp9@1631_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1630 N_OUT9_Mp9@1630_d N_OUT8_Mp9@1630_g N_VDD_Mp9@1630_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1629 N_OUT9_Mn9@1629_d N_OUT8_Mn9@1629_g N_VSS_Mn9@1629_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1628 N_OUT9_Mn9@1628_d N_OUT8_Mn9@1628_g N_VSS_Mn9@1628_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1629 N_OUT9_Mp9@1629_d N_OUT8_Mp9@1629_g N_VDD_Mp9@1629_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1628 N_OUT9_Mp9@1628_d N_OUT8_Mp9@1628_g N_VDD_Mp9@1628_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1627 N_OUT9_Mn9@1627_d N_OUT8_Mn9@1627_g N_VSS_Mn9@1627_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1626 N_OUT9_Mn9@1626_d N_OUT8_Mn9@1626_g N_VSS_Mn9@1626_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1627 N_OUT9_Mp9@1627_d N_OUT8_Mp9@1627_g N_VDD_Mp9@1627_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1626 N_OUT9_Mp9@1626_d N_OUT8_Mp9@1626_g N_VDD_Mp9@1626_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1625 N_OUT9_Mn9@1625_d N_OUT8_Mn9@1625_g N_VSS_Mn9@1625_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1624 N_OUT9_Mn9@1624_d N_OUT8_Mn9@1624_g N_VSS_Mn9@1624_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1625 N_OUT9_Mp9@1625_d N_OUT8_Mp9@1625_g N_VDD_Mp9@1625_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1624 N_OUT9_Mp9@1624_d N_OUT8_Mp9@1624_g N_VDD_Mp9@1624_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1623 N_OUT9_Mn9@1623_d N_OUT8_Mn9@1623_g N_VSS_Mn9@1623_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1622 N_OUT9_Mn9@1622_d N_OUT8_Mn9@1622_g N_VSS_Mn9@1622_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1623 N_OUT9_Mp9@1623_d N_OUT8_Mp9@1623_g N_VDD_Mp9@1623_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1622 N_OUT9_Mp9@1622_d N_OUT8_Mp9@1622_g N_VDD_Mp9@1622_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1621 N_OUT9_Mn9@1621_d N_OUT8_Mn9@1621_g N_VSS_Mn9@1621_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1620 N_OUT9_Mn9@1620_d N_OUT8_Mn9@1620_g N_VSS_Mn9@1620_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1621 N_OUT9_Mp9@1621_d N_OUT8_Mp9@1621_g N_VDD_Mp9@1621_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1620 N_OUT9_Mp9@1620_d N_OUT8_Mp9@1620_g N_VDD_Mp9@1620_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1619 N_OUT9_Mn9@1619_d N_OUT8_Mn9@1619_g N_VSS_Mn9@1619_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1618 N_OUT9_Mn9@1618_d N_OUT8_Mn9@1618_g N_VSS_Mn9@1618_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1619 N_OUT9_Mp9@1619_d N_OUT8_Mp9@1619_g N_VDD_Mp9@1619_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1618 N_OUT9_Mp9@1618_d N_OUT8_Mp9@1618_g N_VDD_Mp9@1618_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1617 N_OUT9_Mn9@1617_d N_OUT8_Mn9@1617_g N_VSS_Mn9@1617_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1616 N_OUT9_Mn9@1616_d N_OUT8_Mn9@1616_g N_VSS_Mn9@1616_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1617 N_OUT9_Mp9@1617_d N_OUT8_Mp9@1617_g N_VDD_Mp9@1617_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1616 N_OUT9_Mp9@1616_d N_OUT8_Mp9@1616_g N_VDD_Mp9@1616_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1615 N_OUT9_Mn9@1615_d N_OUT8_Mn9@1615_g N_VSS_Mn9@1615_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1614 N_OUT9_Mn9@1614_d N_OUT8_Mn9@1614_g N_VSS_Mn9@1614_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1615 N_OUT9_Mp9@1615_d N_OUT8_Mp9@1615_g N_VDD_Mp9@1615_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1614 N_OUT9_Mp9@1614_d N_OUT8_Mp9@1614_g N_VDD_Mp9@1614_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1613 N_OUT9_Mn9@1613_d N_OUT8_Mn9@1613_g N_VSS_Mn9@1613_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1612 N_OUT9_Mn9@1612_d N_OUT8_Mn9@1612_g N_VSS_Mn9@1612_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1613 N_OUT9_Mp9@1613_d N_OUT8_Mp9@1613_g N_VDD_Mp9@1613_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1612 N_OUT9_Mp9@1612_d N_OUT8_Mp9@1612_g N_VDD_Mp9@1612_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1611 N_OUT9_Mn9@1611_d N_OUT8_Mn9@1611_g N_VSS_Mn9@1611_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1610 N_OUT9_Mn9@1610_d N_OUT8_Mn9@1610_g N_VSS_Mn9@1610_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1611 N_OUT9_Mp9@1611_d N_OUT8_Mp9@1611_g N_VDD_Mp9@1611_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1610 N_OUT9_Mp9@1610_d N_OUT8_Mp9@1610_g N_VDD_Mp9@1610_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1609 N_OUT9_Mn9@1609_d N_OUT8_Mn9@1609_g N_VSS_Mn9@1609_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1608 N_OUT9_Mn9@1608_d N_OUT8_Mn9@1608_g N_VSS_Mn9@1608_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1609 N_OUT9_Mp9@1609_d N_OUT8_Mp9@1609_g N_VDD_Mp9@1609_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1608 N_OUT9_Mp9@1608_d N_OUT8_Mp9@1608_g N_VDD_Mp9@1608_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1607 N_OUT9_Mn9@1607_d N_OUT8_Mn9@1607_g N_VSS_Mn9@1607_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1606 N_OUT9_Mn9@1606_d N_OUT8_Mn9@1606_g N_VSS_Mn9@1606_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1607 N_OUT9_Mp9@1607_d N_OUT8_Mp9@1607_g N_VDD_Mp9@1607_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1606 N_OUT9_Mp9@1606_d N_OUT8_Mp9@1606_g N_VDD_Mp9@1606_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1605 N_OUT9_Mn9@1605_d N_OUT8_Mn9@1605_g N_VSS_Mn9@1605_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1604 N_OUT9_Mn9@1604_d N_OUT8_Mn9@1604_g N_VSS_Mn9@1604_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1605 N_OUT9_Mp9@1605_d N_OUT8_Mp9@1605_g N_VDD_Mp9@1605_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1604 N_OUT9_Mp9@1604_d N_OUT8_Mp9@1604_g N_VDD_Mp9@1604_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1603 N_OUT9_Mn9@1603_d N_OUT8_Mn9@1603_g N_VSS_Mn9@1603_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1602 N_OUT9_Mn9@1602_d N_OUT8_Mn9@1602_g N_VSS_Mn9@1602_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1603 N_OUT9_Mp9@1603_d N_OUT8_Mp9@1603_g N_VDD_Mp9@1603_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1602 N_OUT9_Mp9@1602_d N_OUT8_Mp9@1602_g N_VDD_Mp9@1602_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1601 N_OUT9_Mn9@1601_d N_OUT8_Mn9@1601_g N_VSS_Mn9@1601_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1600 N_OUT9_Mn9@1600_d N_OUT8_Mn9@1600_g N_VSS_Mn9@1600_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1601 N_OUT9_Mp9@1601_d N_OUT8_Mp9@1601_g N_VDD_Mp9@1601_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1600 N_OUT9_Mp9@1600_d N_OUT8_Mp9@1600_g N_VDD_Mp9@1600_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1599 N_OUT9_Mn9@1599_d N_OUT8_Mn9@1599_g N_VSS_Mn9@1599_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1598 N_OUT9_Mn9@1598_d N_OUT8_Mn9@1598_g N_VSS_Mn9@1598_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1599 N_OUT9_Mp9@1599_d N_OUT8_Mp9@1599_g N_VDD_Mp9@1599_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1598 N_OUT9_Mp9@1598_d N_OUT8_Mp9@1598_g N_VDD_Mp9@1598_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1597 N_OUT9_Mn9@1597_d N_OUT8_Mn9@1597_g N_VSS_Mn9@1597_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1596 N_OUT9_Mn9@1596_d N_OUT8_Mn9@1596_g N_VSS_Mn9@1596_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1597 N_OUT9_Mp9@1597_d N_OUT8_Mp9@1597_g N_VDD_Mp9@1597_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1596 N_OUT9_Mp9@1596_d N_OUT8_Mp9@1596_g N_VDD_Mp9@1596_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1595 N_OUT9_Mn9@1595_d N_OUT8_Mn9@1595_g N_VSS_Mn9@1595_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1594 N_OUT9_Mn9@1594_d N_OUT8_Mn9@1594_g N_VSS_Mn9@1594_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1595 N_OUT9_Mp9@1595_d N_OUT8_Mp9@1595_g N_VDD_Mp9@1595_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1594 N_OUT9_Mp9@1594_d N_OUT8_Mp9@1594_g N_VDD_Mp9@1594_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1593 N_OUT9_Mn9@1593_d N_OUT8_Mn9@1593_g N_VSS_Mn9@1593_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1592 N_OUT9_Mn9@1592_d N_OUT8_Mn9@1592_g N_VSS_Mn9@1592_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1593 N_OUT9_Mp9@1593_d N_OUT8_Mp9@1593_g N_VDD_Mp9@1593_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1592 N_OUT9_Mp9@1592_d N_OUT8_Mp9@1592_g N_VDD_Mp9@1592_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1591 N_OUT9_Mn9@1591_d N_OUT8_Mn9@1591_g N_VSS_Mn9@1591_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1590 N_OUT9_Mn9@1590_d N_OUT8_Mn9@1590_g N_VSS_Mn9@1590_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1591 N_OUT9_Mp9@1591_d N_OUT8_Mp9@1591_g N_VDD_Mp9@1591_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1590 N_OUT9_Mp9@1590_d N_OUT8_Mp9@1590_g N_VDD_Mp9@1590_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1589 N_OUT9_Mn9@1589_d N_OUT8_Mn9@1589_g N_VSS_Mn9@1589_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1588 N_OUT9_Mn9@1588_d N_OUT8_Mn9@1588_g N_VSS_Mn9@1588_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1589 N_OUT9_Mp9@1589_d N_OUT8_Mp9@1589_g N_VDD_Mp9@1589_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1588 N_OUT9_Mp9@1588_d N_OUT8_Mp9@1588_g N_VDD_Mp9@1588_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1587 N_OUT9_Mn9@1587_d N_OUT8_Mn9@1587_g N_VSS_Mn9@1587_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1586 N_OUT9_Mn9@1586_d N_OUT8_Mn9@1586_g N_VSS_Mn9@1586_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1587 N_OUT9_Mp9@1587_d N_OUT8_Mp9@1587_g N_VDD_Mp9@1587_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1586 N_OUT9_Mp9@1586_d N_OUT8_Mp9@1586_g N_VDD_Mp9@1586_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1585 N_OUT9_Mn9@1585_d N_OUT8_Mn9@1585_g N_VSS_Mn9@1585_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1584 N_OUT9_Mn9@1584_d N_OUT8_Mn9@1584_g N_VSS_Mn9@1584_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1585 N_OUT9_Mp9@1585_d N_OUT8_Mp9@1585_g N_VDD_Mp9@1585_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1584 N_OUT9_Mp9@1584_d N_OUT8_Mp9@1584_g N_VDD_Mp9@1584_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1583 N_OUT9_Mn9@1583_d N_OUT8_Mn9@1583_g N_VSS_Mn9@1583_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1582 N_OUT9_Mn9@1582_d N_OUT8_Mn9@1582_g N_VSS_Mn9@1582_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1583 N_OUT9_Mp9@1583_d N_OUT8_Mp9@1583_g N_VDD_Mp9@1583_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1582 N_OUT9_Mp9@1582_d N_OUT8_Mp9@1582_g N_VDD_Mp9@1582_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1581 N_OUT9_Mn9@1581_d N_OUT8_Mn9@1581_g N_VSS_Mn9@1581_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1580 N_OUT9_Mn9@1580_d N_OUT8_Mn9@1580_g N_VSS_Mn9@1580_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1581 N_OUT9_Mp9@1581_d N_OUT8_Mp9@1581_g N_VDD_Mp9@1581_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1580 N_OUT9_Mp9@1580_d N_OUT8_Mp9@1580_g N_VDD_Mp9@1580_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1579 N_OUT9_Mn9@1579_d N_OUT8_Mn9@1579_g N_VSS_Mn9@1579_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1578 N_OUT9_Mn9@1578_d N_OUT8_Mn9@1578_g N_VSS_Mn9@1578_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1579 N_OUT9_Mp9@1579_d N_OUT8_Mp9@1579_g N_VDD_Mp9@1579_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1578 N_OUT9_Mp9@1578_d N_OUT8_Mp9@1578_g N_VDD_Mp9@1578_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1577 N_OUT9_Mn9@1577_d N_OUT8_Mn9@1577_g N_VSS_Mn9@1577_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1576 N_OUT9_Mn9@1576_d N_OUT8_Mn9@1576_g N_VSS_Mn9@1576_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1577 N_OUT9_Mp9@1577_d N_OUT8_Mp9@1577_g N_VDD_Mp9@1577_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1576 N_OUT9_Mp9@1576_d N_OUT8_Mp9@1576_g N_VDD_Mp9@1576_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1575 N_OUT9_Mn9@1575_d N_OUT8_Mn9@1575_g N_VSS_Mn9@1575_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1574 N_OUT9_Mn9@1574_d N_OUT8_Mn9@1574_g N_VSS_Mn9@1574_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1575 N_OUT9_Mp9@1575_d N_OUT8_Mp9@1575_g N_VDD_Mp9@1575_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1574 N_OUT9_Mp9@1574_d N_OUT8_Mp9@1574_g N_VDD_Mp9@1574_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1573 N_OUT9_Mn9@1573_d N_OUT8_Mn9@1573_g N_VSS_Mn9@1573_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1572 N_OUT9_Mn9@1572_d N_OUT8_Mn9@1572_g N_VSS_Mn9@1572_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1573 N_OUT9_Mp9@1573_d N_OUT8_Mp9@1573_g N_VDD_Mp9@1573_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1572 N_OUT9_Mp9@1572_d N_OUT8_Mp9@1572_g N_VDD_Mp9@1572_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1571 N_OUT9_Mn9@1571_d N_OUT8_Mn9@1571_g N_VSS_Mn9@1571_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1570 N_OUT9_Mn9@1570_d N_OUT8_Mn9@1570_g N_VSS_Mn9@1570_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1571 N_OUT9_Mp9@1571_d N_OUT8_Mp9@1571_g N_VDD_Mp9@1571_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1570 N_OUT9_Mp9@1570_d N_OUT8_Mp9@1570_g N_VDD_Mp9@1570_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1569 N_OUT9_Mn9@1569_d N_OUT8_Mn9@1569_g N_VSS_Mn9@1569_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1568 N_OUT9_Mn9@1568_d N_OUT8_Mn9@1568_g N_VSS_Mn9@1568_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1569 N_OUT9_Mp9@1569_d N_OUT8_Mp9@1569_g N_VDD_Mp9@1569_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1568 N_OUT9_Mp9@1568_d N_OUT8_Mp9@1568_g N_VDD_Mp9@1568_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1567 N_OUT9_Mn9@1567_d N_OUT8_Mn9@1567_g N_VSS_Mn9@1567_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1566 N_OUT9_Mn9@1566_d N_OUT8_Mn9@1566_g N_VSS_Mn9@1566_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1567 N_OUT9_Mp9@1567_d N_OUT8_Mp9@1567_g N_VDD_Mp9@1567_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1566 N_OUT9_Mp9@1566_d N_OUT8_Mp9@1566_g N_VDD_Mp9@1566_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1565 N_OUT9_Mn9@1565_d N_OUT8_Mn9@1565_g N_VSS_Mn9@1565_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1564 N_OUT9_Mn9@1564_d N_OUT8_Mn9@1564_g N_VSS_Mn9@1564_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1565 N_OUT9_Mp9@1565_d N_OUT8_Mp9@1565_g N_VDD_Mp9@1565_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1564 N_OUT9_Mp9@1564_d N_OUT8_Mp9@1564_g N_VDD_Mp9@1564_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1563 N_OUT9_Mn9@1563_d N_OUT8_Mn9@1563_g N_VSS_Mn9@1563_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1562 N_OUT9_Mn9@1562_d N_OUT8_Mn9@1562_g N_VSS_Mn9@1562_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1563 N_OUT9_Mp9@1563_d N_OUT8_Mp9@1563_g N_VDD_Mp9@1563_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1562 N_OUT9_Mp9@1562_d N_OUT8_Mp9@1562_g N_VDD_Mp9@1562_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1561 N_OUT9_Mn9@1561_d N_OUT8_Mn9@1561_g N_VSS_Mn9@1561_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1560 N_OUT9_Mn9@1560_d N_OUT8_Mn9@1560_g N_VSS_Mn9@1560_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1561 N_OUT9_Mp9@1561_d N_OUT8_Mp9@1561_g N_VDD_Mp9@1561_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1560 N_OUT9_Mp9@1560_d N_OUT8_Mp9@1560_g N_VDD_Mp9@1560_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1559 N_OUT9_Mn9@1559_d N_OUT8_Mn9@1559_g N_VSS_Mn9@1559_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1558 N_OUT9_Mn9@1558_d N_OUT8_Mn9@1558_g N_VSS_Mn9@1558_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1559 N_OUT9_Mp9@1559_d N_OUT8_Mp9@1559_g N_VDD_Mp9@1559_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1558 N_OUT9_Mp9@1558_d N_OUT8_Mp9@1558_g N_VDD_Mp9@1558_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1557 N_OUT9_Mn9@1557_d N_OUT8_Mn9@1557_g N_VSS_Mn9@1557_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1556 N_OUT9_Mn9@1556_d N_OUT8_Mn9@1556_g N_VSS_Mn9@1556_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1557 N_OUT9_Mp9@1557_d N_OUT8_Mp9@1557_g N_VDD_Mp9@1557_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1556 N_OUT9_Mp9@1556_d N_OUT8_Mp9@1556_g N_VDD_Mp9@1556_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1555 N_OUT9_Mn9@1555_d N_OUT8_Mn9@1555_g N_VSS_Mn9@1555_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1554 N_OUT9_Mn9@1554_d N_OUT8_Mn9@1554_g N_VSS_Mn9@1554_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1555 N_OUT9_Mp9@1555_d N_OUT8_Mp9@1555_g N_VDD_Mp9@1555_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1554 N_OUT9_Mp9@1554_d N_OUT8_Mp9@1554_g N_VDD_Mp9@1554_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1553 N_OUT9_Mn9@1553_d N_OUT8_Mn9@1553_g N_VSS_Mn9@1553_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1552 N_OUT9_Mn9@1552_d N_OUT8_Mn9@1552_g N_VSS_Mn9@1552_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1553 N_OUT9_Mp9@1553_d N_OUT8_Mp9@1553_g N_VDD_Mp9@1553_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1552 N_OUT9_Mp9@1552_d N_OUT8_Mp9@1552_g N_VDD_Mp9@1552_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1551 N_OUT9_Mn9@1551_d N_OUT8_Mn9@1551_g N_VSS_Mn9@1551_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1550 N_OUT9_Mn9@1550_d N_OUT8_Mn9@1550_g N_VSS_Mn9@1550_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1551 N_OUT9_Mp9@1551_d N_OUT8_Mp9@1551_g N_VDD_Mp9@1551_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1550 N_OUT9_Mp9@1550_d N_OUT8_Mp9@1550_g N_VDD_Mp9@1550_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1549 N_OUT9_Mn9@1549_d N_OUT8_Mn9@1549_g N_VSS_Mn9@1549_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1548 N_OUT9_Mn9@1548_d N_OUT8_Mn9@1548_g N_VSS_Mn9@1548_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1549 N_OUT9_Mp9@1549_d N_OUT8_Mp9@1549_g N_VDD_Mp9@1549_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1548 N_OUT9_Mp9@1548_d N_OUT8_Mp9@1548_g N_VDD_Mp9@1548_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1547 N_OUT9_Mn9@1547_d N_OUT8_Mn9@1547_g N_VSS_Mn9@1547_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1546 N_OUT9_Mn9@1546_d N_OUT8_Mn9@1546_g N_VSS_Mn9@1546_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1547 N_OUT9_Mp9@1547_d N_OUT8_Mp9@1547_g N_VDD_Mp9@1547_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1546 N_OUT9_Mp9@1546_d N_OUT8_Mp9@1546_g N_VDD_Mp9@1546_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1545 N_OUT9_Mn9@1545_d N_OUT8_Mn9@1545_g N_VSS_Mn9@1545_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1544 N_OUT9_Mn9@1544_d N_OUT8_Mn9@1544_g N_VSS_Mn9@1544_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1545 N_OUT9_Mp9@1545_d N_OUT8_Mp9@1545_g N_VDD_Mp9@1545_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1544 N_OUT9_Mp9@1544_d N_OUT8_Mp9@1544_g N_VDD_Mp9@1544_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1543 N_OUT9_Mn9@1543_d N_OUT8_Mn9@1543_g N_VSS_Mn9@1543_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1542 N_OUT9_Mn9@1542_d N_OUT8_Mn9@1542_g N_VSS_Mn9@1542_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1543 N_OUT9_Mp9@1543_d N_OUT8_Mp9@1543_g N_VDD_Mp9@1543_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1542 N_OUT9_Mp9@1542_d N_OUT8_Mp9@1542_g N_VDD_Mp9@1542_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1541 N_OUT9_Mn9@1541_d N_OUT8_Mn9@1541_g N_VSS_Mn9@1541_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1540 N_OUT9_Mn9@1540_d N_OUT8_Mn9@1540_g N_VSS_Mn9@1540_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1541 N_OUT9_Mp9@1541_d N_OUT8_Mp9@1541_g N_VDD_Mp9@1541_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1540 N_OUT9_Mp9@1540_d N_OUT8_Mp9@1540_g N_VDD_Mp9@1540_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1539 N_OUT9_Mn9@1539_d N_OUT8_Mn9@1539_g N_VSS_Mn9@1539_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1538 N_OUT9_Mn9@1538_d N_OUT8_Mn9@1538_g N_VSS_Mn9@1538_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1539 N_OUT9_Mp9@1539_d N_OUT8_Mp9@1539_g N_VDD_Mp9@1539_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1538 N_OUT9_Mp9@1538_d N_OUT8_Mp9@1538_g N_VDD_Mp9@1538_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1537 N_OUT9_Mn9@1537_d N_OUT8_Mn9@1537_g N_VSS_Mn9@1537_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1536 N_OUT9_Mn9@1536_d N_OUT8_Mn9@1536_g N_VSS_Mn9@1536_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1537 N_OUT9_Mp9@1537_d N_OUT8_Mp9@1537_g N_VDD_Mp9@1537_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1536 N_OUT9_Mp9@1536_d N_OUT8_Mp9@1536_g N_VDD_Mp9@1536_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1535 N_OUT9_Mn9@1535_d N_OUT8_Mn9@1535_g N_VSS_Mn9@1535_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1534 N_OUT9_Mn9@1534_d N_OUT8_Mn9@1534_g N_VSS_Mn9@1534_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1535 N_OUT9_Mp9@1535_d N_OUT8_Mp9@1535_g N_VDD_Mp9@1535_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1534 N_OUT9_Mp9@1534_d N_OUT8_Mp9@1534_g N_VDD_Mp9@1534_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1533 N_OUT9_Mn9@1533_d N_OUT8_Mn9@1533_g N_VSS_Mn9@1533_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1532 N_OUT9_Mn9@1532_d N_OUT8_Mn9@1532_g N_VSS_Mn9@1532_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1533 N_OUT9_Mp9@1533_d N_OUT8_Mp9@1533_g N_VDD_Mp9@1533_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1532 N_OUT9_Mp9@1532_d N_OUT8_Mp9@1532_g N_VDD_Mp9@1532_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1531 N_OUT9_Mn9@1531_d N_OUT8_Mn9@1531_g N_VSS_Mn9@1531_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1530 N_OUT9_Mn9@1530_d N_OUT8_Mn9@1530_g N_VSS_Mn9@1530_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1531 N_OUT9_Mp9@1531_d N_OUT8_Mp9@1531_g N_VDD_Mp9@1531_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1530 N_OUT9_Mp9@1530_d N_OUT8_Mp9@1530_g N_VDD_Mp9@1530_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1529 N_OUT9_Mn9@1529_d N_OUT8_Mn9@1529_g N_VSS_Mn9@1529_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1528 N_OUT9_Mn9@1528_d N_OUT8_Mn9@1528_g N_VSS_Mn9@1528_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1529 N_OUT9_Mp9@1529_d N_OUT8_Mp9@1529_g N_VDD_Mp9@1529_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1528 N_OUT9_Mp9@1528_d N_OUT8_Mp9@1528_g N_VDD_Mp9@1528_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1527 N_OUT9_Mn9@1527_d N_OUT8_Mn9@1527_g N_VSS_Mn9@1527_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1526 N_OUT9_Mn9@1526_d N_OUT8_Mn9@1526_g N_VSS_Mn9@1526_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1527 N_OUT9_Mp9@1527_d N_OUT8_Mp9@1527_g N_VDD_Mp9@1527_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1526 N_OUT9_Mp9@1526_d N_OUT8_Mp9@1526_g N_VDD_Mp9@1526_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1525 N_OUT9_Mn9@1525_d N_OUT8_Mn9@1525_g N_VSS_Mn9@1525_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1524 N_OUT9_Mn9@1524_d N_OUT8_Mn9@1524_g N_VSS_Mn9@1524_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1525 N_OUT9_Mp9@1525_d N_OUT8_Mp9@1525_g N_VDD_Mp9@1525_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1524 N_OUT9_Mp9@1524_d N_OUT8_Mp9@1524_g N_VDD_Mp9@1524_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1523 N_OUT9_Mn9@1523_d N_OUT8_Mn9@1523_g N_VSS_Mn9@1523_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1522 N_OUT9_Mn9@1522_d N_OUT8_Mn9@1522_g N_VSS_Mn9@1522_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1523 N_OUT9_Mp9@1523_d N_OUT8_Mp9@1523_g N_VDD_Mp9@1523_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1522 N_OUT9_Mp9@1522_d N_OUT8_Mp9@1522_g N_VDD_Mp9@1522_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1521 N_OUT9_Mn9@1521_d N_OUT8_Mn9@1521_g N_VSS_Mn9@1521_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1520 N_OUT9_Mn9@1520_d N_OUT8_Mn9@1520_g N_VSS_Mn9@1520_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1521 N_OUT9_Mp9@1521_d N_OUT8_Mp9@1521_g N_VDD_Mp9@1521_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1520 N_OUT9_Mp9@1520_d N_OUT8_Mp9@1520_g N_VDD_Mp9@1520_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1519 N_OUT9_Mn9@1519_d N_OUT8_Mn9@1519_g N_VSS_Mn9@1519_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1518 N_OUT9_Mn9@1518_d N_OUT8_Mn9@1518_g N_VSS_Mn9@1518_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1519 N_OUT9_Mp9@1519_d N_OUT8_Mp9@1519_g N_VDD_Mp9@1519_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1518 N_OUT9_Mp9@1518_d N_OUT8_Mp9@1518_g N_VDD_Mp9@1518_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1517 N_OUT9_Mn9@1517_d N_OUT8_Mn9@1517_g N_VSS_Mn9@1517_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1516 N_OUT9_Mn9@1516_d N_OUT8_Mn9@1516_g N_VSS_Mn9@1516_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1517 N_OUT9_Mp9@1517_d N_OUT8_Mp9@1517_g N_VDD_Mp9@1517_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1516 N_OUT9_Mp9@1516_d N_OUT8_Mp9@1516_g N_VDD_Mp9@1516_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1515 N_OUT9_Mn9@1515_d N_OUT8_Mn9@1515_g N_VSS_Mn9@1515_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1514 N_OUT9_Mn9@1514_d N_OUT8_Mn9@1514_g N_VSS_Mn9@1514_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1515 N_OUT9_Mp9@1515_d N_OUT8_Mp9@1515_g N_VDD_Mp9@1515_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1514 N_OUT9_Mp9@1514_d N_OUT8_Mp9@1514_g N_VDD_Mp9@1514_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1513 N_OUT9_Mn9@1513_d N_OUT8_Mn9@1513_g N_VSS_Mn9@1513_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1512 N_OUT9_Mn9@1512_d N_OUT8_Mn9@1512_g N_VSS_Mn9@1512_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1513 N_OUT9_Mp9@1513_d N_OUT8_Mp9@1513_g N_VDD_Mp9@1513_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1512 N_OUT9_Mp9@1512_d N_OUT8_Mp9@1512_g N_VDD_Mp9@1512_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1511 N_OUT9_Mn9@1511_d N_OUT8_Mn9@1511_g N_VSS_Mn9@1511_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1510 N_OUT9_Mn9@1510_d N_OUT8_Mn9@1510_g N_VSS_Mn9@1510_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1511 N_OUT9_Mp9@1511_d N_OUT8_Mp9@1511_g N_VDD_Mp9@1511_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1510 N_OUT9_Mp9@1510_d N_OUT8_Mp9@1510_g N_VDD_Mp9@1510_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1509 N_OUT9_Mn9@1509_d N_OUT8_Mn9@1509_g N_VSS_Mn9@1509_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1508 N_OUT9_Mn9@1508_d N_OUT8_Mn9@1508_g N_VSS_Mn9@1508_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1509 N_OUT9_Mp9@1509_d N_OUT8_Mp9@1509_g N_VDD_Mp9@1509_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1508 N_OUT9_Mp9@1508_d N_OUT8_Mp9@1508_g N_VDD_Mp9@1508_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1507 N_OUT9_Mn9@1507_d N_OUT8_Mn9@1507_g N_VSS_Mn9@1507_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1506 N_OUT9_Mn9@1506_d N_OUT8_Mn9@1506_g N_VSS_Mn9@1506_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1507 N_OUT9_Mp9@1507_d N_OUT8_Mp9@1507_g N_VDD_Mp9@1507_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1506 N_OUT9_Mp9@1506_d N_OUT8_Mp9@1506_g N_VDD_Mp9@1506_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1505 N_OUT9_Mn9@1505_d N_OUT8_Mn9@1505_g N_VSS_Mn9@1505_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1504 N_OUT9_Mn9@1504_d N_OUT8_Mn9@1504_g N_VSS_Mn9@1504_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1505 N_OUT9_Mp9@1505_d N_OUT8_Mp9@1505_g N_VDD_Mp9@1505_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1504 N_OUT9_Mp9@1504_d N_OUT8_Mp9@1504_g N_VDD_Mp9@1504_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1503 N_OUT9_Mn9@1503_d N_OUT8_Mn9@1503_g N_VSS_Mn9@1503_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1502 N_OUT9_Mn9@1502_d N_OUT8_Mn9@1502_g N_VSS_Mn9@1502_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1503 N_OUT9_Mp9@1503_d N_OUT8_Mp9@1503_g N_VDD_Mp9@1503_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1502 N_OUT9_Mp9@1502_d N_OUT8_Mp9@1502_g N_VDD_Mp9@1502_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1501 N_OUT9_Mn9@1501_d N_OUT8_Mn9@1501_g N_VSS_Mn9@1501_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1500 N_OUT9_Mn9@1500_d N_OUT8_Mn9@1500_g N_VSS_Mn9@1500_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1501 N_OUT9_Mp9@1501_d N_OUT8_Mp9@1501_g N_VDD_Mp9@1501_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1500 N_OUT9_Mp9@1500_d N_OUT8_Mp9@1500_g N_VDD_Mp9@1500_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1499 N_OUT9_Mn9@1499_d N_OUT8_Mn9@1499_g N_VSS_Mn9@1499_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1498 N_OUT9_Mn9@1498_d N_OUT8_Mn9@1498_g N_VSS_Mn9@1498_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1499 N_OUT9_Mp9@1499_d N_OUT8_Mp9@1499_g N_VDD_Mp9@1499_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1498 N_OUT9_Mp9@1498_d N_OUT8_Mp9@1498_g N_VDD_Mp9@1498_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1497 N_OUT9_Mn9@1497_d N_OUT8_Mn9@1497_g N_VSS_Mn9@1497_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1496 N_OUT9_Mn9@1496_d N_OUT8_Mn9@1496_g N_VSS_Mn9@1496_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1497 N_OUT9_Mp9@1497_d N_OUT8_Mp9@1497_g N_VDD_Mp9@1497_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1496 N_OUT9_Mp9@1496_d N_OUT8_Mp9@1496_g N_VDD_Mp9@1496_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1495 N_OUT9_Mn9@1495_d N_OUT8_Mn9@1495_g N_VSS_Mn9@1495_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1494 N_OUT9_Mn9@1494_d N_OUT8_Mn9@1494_g N_VSS_Mn9@1494_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1495 N_OUT9_Mp9@1495_d N_OUT8_Mp9@1495_g N_VDD_Mp9@1495_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1494 N_OUT9_Mp9@1494_d N_OUT8_Mp9@1494_g N_VDD_Mp9@1494_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1493 N_OUT9_Mn9@1493_d N_OUT8_Mn9@1493_g N_VSS_Mn9@1493_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1492 N_OUT9_Mn9@1492_d N_OUT8_Mn9@1492_g N_VSS_Mn9@1492_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1493 N_OUT9_Mp9@1493_d N_OUT8_Mp9@1493_g N_VDD_Mp9@1493_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1492 N_OUT9_Mp9@1492_d N_OUT8_Mp9@1492_g N_VDD_Mp9@1492_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1491 N_OUT9_Mn9@1491_d N_OUT8_Mn9@1491_g N_VSS_Mn9@1491_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1490 N_OUT9_Mn9@1490_d N_OUT8_Mn9@1490_g N_VSS_Mn9@1490_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1491 N_OUT9_Mp9@1491_d N_OUT8_Mp9@1491_g N_VDD_Mp9@1491_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1490 N_OUT9_Mp9@1490_d N_OUT8_Mp9@1490_g N_VDD_Mp9@1490_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1489 N_OUT9_Mn9@1489_d N_OUT8_Mn9@1489_g N_VSS_Mn9@1489_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1488 N_OUT9_Mn9@1488_d N_OUT8_Mn9@1488_g N_VSS_Mn9@1488_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1489 N_OUT9_Mp9@1489_d N_OUT8_Mp9@1489_g N_VDD_Mp9@1489_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1488 N_OUT9_Mp9@1488_d N_OUT8_Mp9@1488_g N_VDD_Mp9@1488_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1487 N_OUT9_Mn9@1487_d N_OUT8_Mn9@1487_g N_VSS_Mn9@1487_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1486 N_OUT9_Mn9@1486_d N_OUT8_Mn9@1486_g N_VSS_Mn9@1486_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1487 N_OUT9_Mp9@1487_d N_OUT8_Mp9@1487_g N_VDD_Mp9@1487_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1486 N_OUT9_Mp9@1486_d N_OUT8_Mp9@1486_g N_VDD_Mp9@1486_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1485 N_OUT9_Mn9@1485_d N_OUT8_Mn9@1485_g N_VSS_Mn9@1485_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1484 N_OUT9_Mn9@1484_d N_OUT8_Mn9@1484_g N_VSS_Mn9@1484_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1485 N_OUT9_Mp9@1485_d N_OUT8_Mp9@1485_g N_VDD_Mp9@1485_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1484 N_OUT9_Mp9@1484_d N_OUT8_Mp9@1484_g N_VDD_Mp9@1484_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1483 N_OUT9_Mn9@1483_d N_OUT8_Mn9@1483_g N_VSS_Mn9@1483_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1482 N_OUT9_Mn9@1482_d N_OUT8_Mn9@1482_g N_VSS_Mn9@1482_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1483 N_OUT9_Mp9@1483_d N_OUT8_Mp9@1483_g N_VDD_Mp9@1483_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1482 N_OUT9_Mp9@1482_d N_OUT8_Mp9@1482_g N_VDD_Mp9@1482_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1481 N_OUT9_Mn9@1481_d N_OUT8_Mn9@1481_g N_VSS_Mn9@1481_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1480 N_OUT9_Mn9@1480_d N_OUT8_Mn9@1480_g N_VSS_Mn9@1480_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1481 N_OUT9_Mp9@1481_d N_OUT8_Mp9@1481_g N_VDD_Mp9@1481_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1480 N_OUT9_Mp9@1480_d N_OUT8_Mp9@1480_g N_VDD_Mp9@1480_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1479 N_OUT9_Mn9@1479_d N_OUT8_Mn9@1479_g N_VSS_Mn9@1479_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1478 N_OUT9_Mn9@1478_d N_OUT8_Mn9@1478_g N_VSS_Mn9@1478_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1479 N_OUT9_Mp9@1479_d N_OUT8_Mp9@1479_g N_VDD_Mp9@1479_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1478 N_OUT9_Mp9@1478_d N_OUT8_Mp9@1478_g N_VDD_Mp9@1478_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1477 N_OUT9_Mn9@1477_d N_OUT8_Mn9@1477_g N_VSS_Mn9@1477_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1476 N_OUT9_Mn9@1476_d N_OUT8_Mn9@1476_g N_VSS_Mn9@1476_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1477 N_OUT9_Mp9@1477_d N_OUT8_Mp9@1477_g N_VDD_Mp9@1477_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1476 N_OUT9_Mp9@1476_d N_OUT8_Mp9@1476_g N_VDD_Mp9@1476_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1475 N_OUT9_Mn9@1475_d N_OUT8_Mn9@1475_g N_VSS_Mn9@1475_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1474 N_OUT9_Mn9@1474_d N_OUT8_Mn9@1474_g N_VSS_Mn9@1474_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1475 N_OUT9_Mp9@1475_d N_OUT8_Mp9@1475_g N_VDD_Mp9@1475_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1474 N_OUT9_Mp9@1474_d N_OUT8_Mp9@1474_g N_VDD_Mp9@1474_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1473 N_OUT9_Mn9@1473_d N_OUT8_Mn9@1473_g N_VSS_Mn9@1473_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1472 N_OUT9_Mn9@1472_d N_OUT8_Mn9@1472_g N_VSS_Mn9@1472_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1473 N_OUT9_Mp9@1473_d N_OUT8_Mp9@1473_g N_VDD_Mp9@1473_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1472 N_OUT9_Mp9@1472_d N_OUT8_Mp9@1472_g N_VDD_Mp9@1472_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1471 N_OUT9_Mn9@1471_d N_OUT8_Mn9@1471_g N_VSS_Mn9@1471_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1470 N_OUT9_Mn9@1470_d N_OUT8_Mn9@1470_g N_VSS_Mn9@1470_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1471 N_OUT9_Mp9@1471_d N_OUT8_Mp9@1471_g N_VDD_Mp9@1471_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1470 N_OUT9_Mp9@1470_d N_OUT8_Mp9@1470_g N_VDD_Mp9@1470_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1469 N_OUT9_Mn9@1469_d N_OUT8_Mn9@1469_g N_VSS_Mn9@1469_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1468 N_OUT9_Mn9@1468_d N_OUT8_Mn9@1468_g N_VSS_Mn9@1468_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1469 N_OUT9_Mp9@1469_d N_OUT8_Mp9@1469_g N_VDD_Mp9@1469_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1468 N_OUT9_Mp9@1468_d N_OUT8_Mp9@1468_g N_VDD_Mp9@1468_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1467 N_OUT9_Mn9@1467_d N_OUT8_Mn9@1467_g N_VSS_Mn9@1467_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1466 N_OUT9_Mn9@1466_d N_OUT8_Mn9@1466_g N_VSS_Mn9@1466_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1467 N_OUT9_Mp9@1467_d N_OUT8_Mp9@1467_g N_VDD_Mp9@1467_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1466 N_OUT9_Mp9@1466_d N_OUT8_Mp9@1466_g N_VDD_Mp9@1466_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1465 N_OUT9_Mn9@1465_d N_OUT8_Mn9@1465_g N_VSS_Mn9@1465_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1464 N_OUT9_Mn9@1464_d N_OUT8_Mn9@1464_g N_VSS_Mn9@1464_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1465 N_OUT9_Mp9@1465_d N_OUT8_Mp9@1465_g N_VDD_Mp9@1465_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1464 N_OUT9_Mp9@1464_d N_OUT8_Mp9@1464_g N_VDD_Mp9@1464_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1463 N_OUT9_Mn9@1463_d N_OUT8_Mn9@1463_g N_VSS_Mn9@1463_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1462 N_OUT9_Mn9@1462_d N_OUT8_Mn9@1462_g N_VSS_Mn9@1462_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1463 N_OUT9_Mp9@1463_d N_OUT8_Mp9@1463_g N_VDD_Mp9@1463_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1462 N_OUT9_Mp9@1462_d N_OUT8_Mp9@1462_g N_VDD_Mp9@1462_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1461 N_OUT9_Mn9@1461_d N_OUT8_Mn9@1461_g N_VSS_Mn9@1461_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1460 N_OUT9_Mn9@1460_d N_OUT8_Mn9@1460_g N_VSS_Mn9@1460_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1461 N_OUT9_Mp9@1461_d N_OUT8_Mp9@1461_g N_VDD_Mp9@1461_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1460 N_OUT9_Mp9@1460_d N_OUT8_Mp9@1460_g N_VDD_Mp9@1460_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1459 N_OUT9_Mn9@1459_d N_OUT8_Mn9@1459_g N_VSS_Mn9@1459_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1458 N_OUT9_Mn9@1458_d N_OUT8_Mn9@1458_g N_VSS_Mn9@1458_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1459 N_OUT9_Mp9@1459_d N_OUT8_Mp9@1459_g N_VDD_Mp9@1459_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1458 N_OUT9_Mp9@1458_d N_OUT8_Mp9@1458_g N_VDD_Mp9@1458_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1457 N_OUT9_Mn9@1457_d N_OUT8_Mn9@1457_g N_VSS_Mn9@1457_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1456 N_OUT9_Mn9@1456_d N_OUT8_Mn9@1456_g N_VSS_Mn9@1456_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1457 N_OUT9_Mp9@1457_d N_OUT8_Mp9@1457_g N_VDD_Mp9@1457_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1456 N_OUT9_Mp9@1456_d N_OUT8_Mp9@1456_g N_VDD_Mp9@1456_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1455 N_OUT9_Mn9@1455_d N_OUT8_Mn9@1455_g N_VSS_Mn9@1455_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1454 N_OUT9_Mn9@1454_d N_OUT8_Mn9@1454_g N_VSS_Mn9@1454_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1455 N_OUT9_Mp9@1455_d N_OUT8_Mp9@1455_g N_VDD_Mp9@1455_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1454 N_OUT9_Mp9@1454_d N_OUT8_Mp9@1454_g N_VDD_Mp9@1454_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1453 N_OUT9_Mn9@1453_d N_OUT8_Mn9@1453_g N_VSS_Mn9@1453_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1452 N_OUT9_Mn9@1452_d N_OUT8_Mn9@1452_g N_VSS_Mn9@1452_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1453 N_OUT9_Mp9@1453_d N_OUT8_Mp9@1453_g N_VDD_Mp9@1453_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1452 N_OUT9_Mp9@1452_d N_OUT8_Mp9@1452_g N_VDD_Mp9@1452_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1451 N_OUT9_Mn9@1451_d N_OUT8_Mn9@1451_g N_VSS_Mn9@1451_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1450 N_OUT9_Mn9@1450_d N_OUT8_Mn9@1450_g N_VSS_Mn9@1450_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1451 N_OUT9_Mp9@1451_d N_OUT8_Mp9@1451_g N_VDD_Mp9@1451_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1450 N_OUT9_Mp9@1450_d N_OUT8_Mp9@1450_g N_VDD_Mp9@1450_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1449 N_OUT9_Mn9@1449_d N_OUT8_Mn9@1449_g N_VSS_Mn9@1449_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1448 N_OUT9_Mn9@1448_d N_OUT8_Mn9@1448_g N_VSS_Mn9@1448_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1449 N_OUT9_Mp9@1449_d N_OUT8_Mp9@1449_g N_VDD_Mp9@1449_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1448 N_OUT9_Mp9@1448_d N_OUT8_Mp9@1448_g N_VDD_Mp9@1448_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1447 N_OUT9_Mn9@1447_d N_OUT8_Mn9@1447_g N_VSS_Mn9@1447_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1446 N_OUT9_Mn9@1446_d N_OUT8_Mn9@1446_g N_VSS_Mn9@1446_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1447 N_OUT9_Mp9@1447_d N_OUT8_Mp9@1447_g N_VDD_Mp9@1447_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1446 N_OUT9_Mp9@1446_d N_OUT8_Mp9@1446_g N_VDD_Mp9@1446_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1445 N_OUT9_Mn9@1445_d N_OUT8_Mn9@1445_g N_VSS_Mn9@1445_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1444 N_OUT9_Mn9@1444_d N_OUT8_Mn9@1444_g N_VSS_Mn9@1444_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1445 N_OUT9_Mp9@1445_d N_OUT8_Mp9@1445_g N_VDD_Mp9@1445_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1444 N_OUT9_Mp9@1444_d N_OUT8_Mp9@1444_g N_VDD_Mp9@1444_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1443 N_OUT9_Mn9@1443_d N_OUT8_Mn9@1443_g N_VSS_Mn9@1443_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1442 N_OUT9_Mn9@1442_d N_OUT8_Mn9@1442_g N_VSS_Mn9@1442_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1443 N_OUT9_Mp9@1443_d N_OUT8_Mp9@1443_g N_VDD_Mp9@1443_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1442 N_OUT9_Mp9@1442_d N_OUT8_Mp9@1442_g N_VDD_Mp9@1442_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1441 N_OUT9_Mn9@1441_d N_OUT8_Mn9@1441_g N_VSS_Mn9@1441_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1440 N_OUT9_Mn9@1440_d N_OUT8_Mn9@1440_g N_VSS_Mn9@1440_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1441 N_OUT9_Mp9@1441_d N_OUT8_Mp9@1441_g N_VDD_Mp9@1441_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1440 N_OUT9_Mp9@1440_d N_OUT8_Mp9@1440_g N_VDD_Mp9@1440_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1439 N_OUT9_Mn9@1439_d N_OUT8_Mn9@1439_g N_VSS_Mn9@1439_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1438 N_OUT9_Mn9@1438_d N_OUT8_Mn9@1438_g N_VSS_Mn9@1438_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1439 N_OUT9_Mp9@1439_d N_OUT8_Mp9@1439_g N_VDD_Mp9@1439_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1438 N_OUT9_Mp9@1438_d N_OUT8_Mp9@1438_g N_VDD_Mp9@1438_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1437 N_OUT9_Mn9@1437_d N_OUT8_Mn9@1437_g N_VSS_Mn9@1437_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1436 N_OUT9_Mn9@1436_d N_OUT8_Mn9@1436_g N_VSS_Mn9@1436_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1437 N_OUT9_Mp9@1437_d N_OUT8_Mp9@1437_g N_VDD_Mp9@1437_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1436 N_OUT9_Mp9@1436_d N_OUT8_Mp9@1436_g N_VDD_Mp9@1436_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1435 N_OUT9_Mn9@1435_d N_OUT8_Mn9@1435_g N_VSS_Mn9@1435_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1434 N_OUT9_Mn9@1434_d N_OUT8_Mn9@1434_g N_VSS_Mn9@1434_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1435 N_OUT9_Mp9@1435_d N_OUT8_Mp9@1435_g N_VDD_Mp9@1435_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1434 N_OUT9_Mp9@1434_d N_OUT8_Mp9@1434_g N_VDD_Mp9@1434_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1433 N_OUT9_Mn9@1433_d N_OUT8_Mn9@1433_g N_VSS_Mn9@1433_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1432 N_OUT9_Mn9@1432_d N_OUT8_Mn9@1432_g N_VSS_Mn9@1432_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1433 N_OUT9_Mp9@1433_d N_OUT8_Mp9@1433_g N_VDD_Mp9@1433_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1432 N_OUT9_Mp9@1432_d N_OUT8_Mp9@1432_g N_VDD_Mp9@1432_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1431 N_OUT9_Mn9@1431_d N_OUT8_Mn9@1431_g N_VSS_Mn9@1431_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1430 N_OUT9_Mn9@1430_d N_OUT8_Mn9@1430_g N_VSS_Mn9@1430_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1431 N_OUT9_Mp9@1431_d N_OUT8_Mp9@1431_g N_VDD_Mp9@1431_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1430 N_OUT9_Mp9@1430_d N_OUT8_Mp9@1430_g N_VDD_Mp9@1430_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1429 N_OUT9_Mn9@1429_d N_OUT8_Mn9@1429_g N_VSS_Mn9@1429_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1428 N_OUT9_Mn9@1428_d N_OUT8_Mn9@1428_g N_VSS_Mn9@1428_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1429 N_OUT9_Mp9@1429_d N_OUT8_Mp9@1429_g N_VDD_Mp9@1429_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1428 N_OUT9_Mp9@1428_d N_OUT8_Mp9@1428_g N_VDD_Mp9@1428_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1427 N_OUT9_Mn9@1427_d N_OUT8_Mn9@1427_g N_VSS_Mn9@1427_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1426 N_OUT9_Mn9@1426_d N_OUT8_Mn9@1426_g N_VSS_Mn9@1426_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1427 N_OUT9_Mp9@1427_d N_OUT8_Mp9@1427_g N_VDD_Mp9@1427_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1426 N_OUT9_Mp9@1426_d N_OUT8_Mp9@1426_g N_VDD_Mp9@1426_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1425 N_OUT9_Mn9@1425_d N_OUT8_Mn9@1425_g N_VSS_Mn9@1425_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1424 N_OUT9_Mn9@1424_d N_OUT8_Mn9@1424_g N_VSS_Mn9@1424_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1425 N_OUT9_Mp9@1425_d N_OUT8_Mp9@1425_g N_VDD_Mp9@1425_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1424 N_OUT9_Mp9@1424_d N_OUT8_Mp9@1424_g N_VDD_Mp9@1424_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1423 N_OUT9_Mn9@1423_d N_OUT8_Mn9@1423_g N_VSS_Mn9@1423_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1422 N_OUT9_Mn9@1422_d N_OUT8_Mn9@1422_g N_VSS_Mn9@1422_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1423 N_OUT9_Mp9@1423_d N_OUT8_Mp9@1423_g N_VDD_Mp9@1423_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1422 N_OUT9_Mp9@1422_d N_OUT8_Mp9@1422_g N_VDD_Mp9@1422_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1421 N_OUT9_Mn9@1421_d N_OUT8_Mn9@1421_g N_VSS_Mn9@1421_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1420 N_OUT9_Mn9@1420_d N_OUT8_Mn9@1420_g N_VSS_Mn9@1420_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1421 N_OUT9_Mp9@1421_d N_OUT8_Mp9@1421_g N_VDD_Mp9@1421_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1420 N_OUT9_Mp9@1420_d N_OUT8_Mp9@1420_g N_VDD_Mp9@1420_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1419 N_OUT9_Mn9@1419_d N_OUT8_Mn9@1419_g N_VSS_Mn9@1419_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1418 N_OUT9_Mn9@1418_d N_OUT8_Mn9@1418_g N_VSS_Mn9@1418_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1419 N_OUT9_Mp9@1419_d N_OUT8_Mp9@1419_g N_VDD_Mp9@1419_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1418 N_OUT9_Mp9@1418_d N_OUT8_Mp9@1418_g N_VDD_Mp9@1418_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1417 N_OUT9_Mn9@1417_d N_OUT8_Mn9@1417_g N_VSS_Mn9@1417_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1416 N_OUT9_Mn9@1416_d N_OUT8_Mn9@1416_g N_VSS_Mn9@1416_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1417 N_OUT9_Mp9@1417_d N_OUT8_Mp9@1417_g N_VDD_Mp9@1417_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1416 N_OUT9_Mp9@1416_d N_OUT8_Mp9@1416_g N_VDD_Mp9@1416_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1415 N_OUT9_Mn9@1415_d N_OUT8_Mn9@1415_g N_VSS_Mn9@1415_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1414 N_OUT9_Mn9@1414_d N_OUT8_Mn9@1414_g N_VSS_Mn9@1414_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1415 N_OUT9_Mp9@1415_d N_OUT8_Mp9@1415_g N_VDD_Mp9@1415_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1414 N_OUT9_Mp9@1414_d N_OUT8_Mp9@1414_g N_VDD_Mp9@1414_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1413 N_OUT9_Mn9@1413_d N_OUT8_Mn9@1413_g N_VSS_Mn9@1413_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1412 N_OUT9_Mn9@1412_d N_OUT8_Mn9@1412_g N_VSS_Mn9@1412_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1413 N_OUT9_Mp9@1413_d N_OUT8_Mp9@1413_g N_VDD_Mp9@1413_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1412 N_OUT9_Mp9@1412_d N_OUT8_Mp9@1412_g N_VDD_Mp9@1412_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1411 N_OUT9_Mn9@1411_d N_OUT8_Mn9@1411_g N_VSS_Mn9@1411_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1410 N_OUT9_Mn9@1410_d N_OUT8_Mn9@1410_g N_VSS_Mn9@1410_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1411 N_OUT9_Mp9@1411_d N_OUT8_Mp9@1411_g N_VDD_Mp9@1411_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1410 N_OUT9_Mp9@1410_d N_OUT8_Mp9@1410_g N_VDD_Mp9@1410_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1409 N_OUT9_Mn9@1409_d N_OUT8_Mn9@1409_g N_VSS_Mn9@1409_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1408 N_OUT9_Mn9@1408_d N_OUT8_Mn9@1408_g N_VSS_Mn9@1408_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1409 N_OUT9_Mp9@1409_d N_OUT8_Mp9@1409_g N_VDD_Mp9@1409_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1408 N_OUT9_Mp9@1408_d N_OUT8_Mp9@1408_g N_VDD_Mp9@1408_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1407 N_OUT9_Mn9@1407_d N_OUT8_Mn9@1407_g N_VSS_Mn9@1407_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1406 N_OUT9_Mn9@1406_d N_OUT8_Mn9@1406_g N_VSS_Mn9@1406_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1407 N_OUT9_Mp9@1407_d N_OUT8_Mp9@1407_g N_VDD_Mp9@1407_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1406 N_OUT9_Mp9@1406_d N_OUT8_Mp9@1406_g N_VDD_Mp9@1406_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1405 N_OUT9_Mn9@1405_d N_OUT8_Mn9@1405_g N_VSS_Mn9@1405_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1404 N_OUT9_Mn9@1404_d N_OUT8_Mn9@1404_g N_VSS_Mn9@1404_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1405 N_OUT9_Mp9@1405_d N_OUT8_Mp9@1405_g N_VDD_Mp9@1405_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1404 N_OUT9_Mp9@1404_d N_OUT8_Mp9@1404_g N_VDD_Mp9@1404_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1403 N_OUT9_Mn9@1403_d N_OUT8_Mn9@1403_g N_VSS_Mn9@1403_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1402 N_OUT9_Mn9@1402_d N_OUT8_Mn9@1402_g N_VSS_Mn9@1402_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1403 N_OUT9_Mp9@1403_d N_OUT8_Mp9@1403_g N_VDD_Mp9@1403_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1402 N_OUT9_Mp9@1402_d N_OUT8_Mp9@1402_g N_VDD_Mp9@1402_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1401 N_OUT9_Mn9@1401_d N_OUT8_Mn9@1401_g N_VSS_Mn9@1401_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1400 N_OUT9_Mn9@1400_d N_OUT8_Mn9@1400_g N_VSS_Mn9@1400_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1401 N_OUT9_Mp9@1401_d N_OUT8_Mp9@1401_g N_VDD_Mp9@1401_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1400 N_OUT9_Mp9@1400_d N_OUT8_Mp9@1400_g N_VDD_Mp9@1400_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1399 N_OUT9_Mn9@1399_d N_OUT8_Mn9@1399_g N_VSS_Mn9@1399_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1398 N_OUT9_Mn9@1398_d N_OUT8_Mn9@1398_g N_VSS_Mn9@1398_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1399 N_OUT9_Mp9@1399_d N_OUT8_Mp9@1399_g N_VDD_Mp9@1399_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1398 N_OUT9_Mp9@1398_d N_OUT8_Mp9@1398_g N_VDD_Mp9@1398_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1397 N_OUT9_Mn9@1397_d N_OUT8_Mn9@1397_g N_VSS_Mn9@1397_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1396 N_OUT9_Mn9@1396_d N_OUT8_Mn9@1396_g N_VSS_Mn9@1396_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1397 N_OUT9_Mp9@1397_d N_OUT8_Mp9@1397_g N_VDD_Mp9@1397_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1396 N_OUT9_Mp9@1396_d N_OUT8_Mp9@1396_g N_VDD_Mp9@1396_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1395 N_OUT9_Mn9@1395_d N_OUT8_Mn9@1395_g N_VSS_Mn9@1395_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1394 N_OUT9_Mn9@1394_d N_OUT8_Mn9@1394_g N_VSS_Mn9@1394_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1395 N_OUT9_Mp9@1395_d N_OUT8_Mp9@1395_g N_VDD_Mp9@1395_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1394 N_OUT9_Mp9@1394_d N_OUT8_Mp9@1394_g N_VDD_Mp9@1394_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1393 N_OUT9_Mn9@1393_d N_OUT8_Mn9@1393_g N_VSS_Mn9@1393_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1392 N_OUT9_Mn9@1392_d N_OUT8_Mn9@1392_g N_VSS_Mn9@1392_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1393 N_OUT9_Mp9@1393_d N_OUT8_Mp9@1393_g N_VDD_Mp9@1393_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1392 N_OUT9_Mp9@1392_d N_OUT8_Mp9@1392_g N_VDD_Mp9@1392_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1391 N_OUT9_Mn9@1391_d N_OUT8_Mn9@1391_g N_VSS_Mn9@1391_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1390 N_OUT9_Mn9@1390_d N_OUT8_Mn9@1390_g N_VSS_Mn9@1390_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1391 N_OUT9_Mp9@1391_d N_OUT8_Mp9@1391_g N_VDD_Mp9@1391_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1390 N_OUT9_Mp9@1390_d N_OUT8_Mp9@1390_g N_VDD_Mp9@1390_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1389 N_OUT9_Mn9@1389_d N_OUT8_Mn9@1389_g N_VSS_Mn9@1389_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1388 N_OUT9_Mn9@1388_d N_OUT8_Mn9@1388_g N_VSS_Mn9@1388_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1389 N_OUT9_Mp9@1389_d N_OUT8_Mp9@1389_g N_VDD_Mp9@1389_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1388 N_OUT9_Mp9@1388_d N_OUT8_Mp9@1388_g N_VDD_Mp9@1388_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1387 N_OUT9_Mn9@1387_d N_OUT8_Mn9@1387_g N_VSS_Mn9@1387_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1386 N_OUT9_Mn9@1386_d N_OUT8_Mn9@1386_g N_VSS_Mn9@1386_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1387 N_OUT9_Mp9@1387_d N_OUT8_Mp9@1387_g N_VDD_Mp9@1387_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1386 N_OUT9_Mp9@1386_d N_OUT8_Mp9@1386_g N_VDD_Mp9@1386_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1385 N_OUT9_Mn9@1385_d N_OUT8_Mn9@1385_g N_VSS_Mn9@1385_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1384 N_OUT9_Mn9@1384_d N_OUT8_Mn9@1384_g N_VSS_Mn9@1384_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1385 N_OUT9_Mp9@1385_d N_OUT8_Mp9@1385_g N_VDD_Mp9@1385_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1384 N_OUT9_Mp9@1384_d N_OUT8_Mp9@1384_g N_VDD_Mp9@1384_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1383 N_OUT9_Mn9@1383_d N_OUT8_Mn9@1383_g N_VSS_Mn9@1383_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1382 N_OUT9_Mn9@1382_d N_OUT8_Mn9@1382_g N_VSS_Mn9@1382_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1383 N_OUT9_Mp9@1383_d N_OUT8_Mp9@1383_g N_VDD_Mp9@1383_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1382 N_OUT9_Mp9@1382_d N_OUT8_Mp9@1382_g N_VDD_Mp9@1382_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1381 N_OUT9_Mn9@1381_d N_OUT8_Mn9@1381_g N_VSS_Mn9@1381_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1380 N_OUT9_Mn9@1380_d N_OUT8_Mn9@1380_g N_VSS_Mn9@1380_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1381 N_OUT9_Mp9@1381_d N_OUT8_Mp9@1381_g N_VDD_Mp9@1381_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1380 N_OUT9_Mp9@1380_d N_OUT8_Mp9@1380_g N_VDD_Mp9@1380_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1379 N_OUT9_Mn9@1379_d N_OUT8_Mn9@1379_g N_VSS_Mn9@1379_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1378 N_OUT9_Mn9@1378_d N_OUT8_Mn9@1378_g N_VSS_Mn9@1378_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1379 N_OUT9_Mp9@1379_d N_OUT8_Mp9@1379_g N_VDD_Mp9@1379_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1378 N_OUT9_Mp9@1378_d N_OUT8_Mp9@1378_g N_VDD_Mp9@1378_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1377 N_OUT9_Mn9@1377_d N_OUT8_Mn9@1377_g N_VSS_Mn9@1377_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1376 N_OUT9_Mn9@1376_d N_OUT8_Mn9@1376_g N_VSS_Mn9@1376_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1377 N_OUT9_Mp9@1377_d N_OUT8_Mp9@1377_g N_VDD_Mp9@1377_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1376 N_OUT9_Mp9@1376_d N_OUT8_Mp9@1376_g N_VDD_Mp9@1376_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1375 N_OUT9_Mn9@1375_d N_OUT8_Mn9@1375_g N_VSS_Mn9@1375_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1374 N_OUT9_Mn9@1374_d N_OUT8_Mn9@1374_g N_VSS_Mn9@1374_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1375 N_OUT9_Mp9@1375_d N_OUT8_Mp9@1375_g N_VDD_Mp9@1375_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1374 N_OUT9_Mp9@1374_d N_OUT8_Mp9@1374_g N_VDD_Mp9@1374_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1373 N_OUT9_Mn9@1373_d N_OUT8_Mn9@1373_g N_VSS_Mn9@1373_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1372 N_OUT9_Mn9@1372_d N_OUT8_Mn9@1372_g N_VSS_Mn9@1372_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1373 N_OUT9_Mp9@1373_d N_OUT8_Mp9@1373_g N_VDD_Mp9@1373_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1372 N_OUT9_Mp9@1372_d N_OUT8_Mp9@1372_g N_VDD_Mp9@1372_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1371 N_OUT9_Mn9@1371_d N_OUT8_Mn9@1371_g N_VSS_Mn9@1371_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1370 N_OUT9_Mn9@1370_d N_OUT8_Mn9@1370_g N_VSS_Mn9@1370_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1371 N_OUT9_Mp9@1371_d N_OUT8_Mp9@1371_g N_VDD_Mp9@1371_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1370 N_OUT9_Mp9@1370_d N_OUT8_Mp9@1370_g N_VDD_Mp9@1370_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1369 N_OUT9_Mn9@1369_d N_OUT8_Mn9@1369_g N_VSS_Mn9@1369_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1368 N_OUT9_Mn9@1368_d N_OUT8_Mn9@1368_g N_VSS_Mn9@1368_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1369 N_OUT9_Mp9@1369_d N_OUT8_Mp9@1369_g N_VDD_Mp9@1369_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1368 N_OUT9_Mp9@1368_d N_OUT8_Mp9@1368_g N_VDD_Mp9@1368_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1367 N_OUT9_Mn9@1367_d N_OUT8_Mn9@1367_g N_VSS_Mn9@1367_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1366 N_OUT9_Mn9@1366_d N_OUT8_Mn9@1366_g N_VSS_Mn9@1366_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1367 N_OUT9_Mp9@1367_d N_OUT8_Mp9@1367_g N_VDD_Mp9@1367_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1366 N_OUT9_Mp9@1366_d N_OUT8_Mp9@1366_g N_VDD_Mp9@1366_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1365 N_OUT9_Mn9@1365_d N_OUT8_Mn9@1365_g N_VSS_Mn9@1365_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1364 N_OUT9_Mn9@1364_d N_OUT8_Mn9@1364_g N_VSS_Mn9@1364_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1365 N_OUT9_Mp9@1365_d N_OUT8_Mp9@1365_g N_VDD_Mp9@1365_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1364 N_OUT9_Mp9@1364_d N_OUT8_Mp9@1364_g N_VDD_Mp9@1364_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1363 N_OUT9_Mn9@1363_d N_OUT8_Mn9@1363_g N_VSS_Mn9@1363_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1362 N_OUT9_Mn9@1362_d N_OUT8_Mn9@1362_g N_VSS_Mn9@1362_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1363 N_OUT9_Mp9@1363_d N_OUT8_Mp9@1363_g N_VDD_Mp9@1363_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1362 N_OUT9_Mp9@1362_d N_OUT8_Mp9@1362_g N_VDD_Mp9@1362_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1361 N_OUT9_Mn9@1361_d N_OUT8_Mn9@1361_g N_VSS_Mn9@1361_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1360 N_OUT9_Mn9@1360_d N_OUT8_Mn9@1360_g N_VSS_Mn9@1360_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1361 N_OUT9_Mp9@1361_d N_OUT8_Mp9@1361_g N_VDD_Mp9@1361_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1360 N_OUT9_Mp9@1360_d N_OUT8_Mp9@1360_g N_VDD_Mp9@1360_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1359 N_OUT9_Mn9@1359_d N_OUT8_Mn9@1359_g N_VSS_Mn9@1359_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1358 N_OUT9_Mn9@1358_d N_OUT8_Mn9@1358_g N_VSS_Mn9@1358_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1359 N_OUT9_Mp9@1359_d N_OUT8_Mp9@1359_g N_VDD_Mp9@1359_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1358 N_OUT9_Mp9@1358_d N_OUT8_Mp9@1358_g N_VDD_Mp9@1358_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1357 N_OUT9_Mn9@1357_d N_OUT8_Mn9@1357_g N_VSS_Mn9@1357_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1356 N_OUT9_Mn9@1356_d N_OUT8_Mn9@1356_g N_VSS_Mn9@1356_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1357 N_OUT9_Mp9@1357_d N_OUT8_Mp9@1357_g N_VDD_Mp9@1357_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1356 N_OUT9_Mp9@1356_d N_OUT8_Mp9@1356_g N_VDD_Mp9@1356_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1355 N_OUT9_Mn9@1355_d N_OUT8_Mn9@1355_g N_VSS_Mn9@1355_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1354 N_OUT9_Mn9@1354_d N_OUT8_Mn9@1354_g N_VSS_Mn9@1354_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1355 N_OUT9_Mp9@1355_d N_OUT8_Mp9@1355_g N_VDD_Mp9@1355_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1354 N_OUT9_Mp9@1354_d N_OUT8_Mp9@1354_g N_VDD_Mp9@1354_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1353 N_OUT9_Mn9@1353_d N_OUT8_Mn9@1353_g N_VSS_Mn9@1353_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1352 N_OUT9_Mn9@1352_d N_OUT8_Mn9@1352_g N_VSS_Mn9@1352_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1353 N_OUT9_Mp9@1353_d N_OUT8_Mp9@1353_g N_VDD_Mp9@1353_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1352 N_OUT9_Mp9@1352_d N_OUT8_Mp9@1352_g N_VDD_Mp9@1352_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1351 N_OUT9_Mn9@1351_d N_OUT8_Mn9@1351_g N_VSS_Mn9@1351_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1350 N_OUT9_Mn9@1350_d N_OUT8_Mn9@1350_g N_VSS_Mn9@1350_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1351 N_OUT9_Mp9@1351_d N_OUT8_Mp9@1351_g N_VDD_Mp9@1351_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1350 N_OUT9_Mp9@1350_d N_OUT8_Mp9@1350_g N_VDD_Mp9@1350_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1349 N_OUT9_Mn9@1349_d N_OUT8_Mn9@1349_g N_VSS_Mn9@1349_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1348 N_OUT9_Mn9@1348_d N_OUT8_Mn9@1348_g N_VSS_Mn9@1348_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1349 N_OUT9_Mp9@1349_d N_OUT8_Mp9@1349_g N_VDD_Mp9@1349_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1348 N_OUT9_Mp9@1348_d N_OUT8_Mp9@1348_g N_VDD_Mp9@1348_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1347 N_OUT9_Mn9@1347_d N_OUT8_Mn9@1347_g N_VSS_Mn9@1347_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1346 N_OUT9_Mn9@1346_d N_OUT8_Mn9@1346_g N_VSS_Mn9@1346_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1347 N_OUT9_Mp9@1347_d N_OUT8_Mp9@1347_g N_VDD_Mp9@1347_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1346 N_OUT9_Mp9@1346_d N_OUT8_Mp9@1346_g N_VDD_Mp9@1346_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1345 N_OUT9_Mn9@1345_d N_OUT8_Mn9@1345_g N_VSS_Mn9@1345_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1344 N_OUT9_Mn9@1344_d N_OUT8_Mn9@1344_g N_VSS_Mn9@1344_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1345 N_OUT9_Mp9@1345_d N_OUT8_Mp9@1345_g N_VDD_Mp9@1345_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1344 N_OUT9_Mp9@1344_d N_OUT8_Mp9@1344_g N_VDD_Mp9@1344_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1343 N_OUT9_Mn9@1343_d N_OUT8_Mn9@1343_g N_VSS_Mn9@1343_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1342 N_OUT9_Mn9@1342_d N_OUT8_Mn9@1342_g N_VSS_Mn9@1342_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1343 N_OUT9_Mp9@1343_d N_OUT8_Mp9@1343_g N_VDD_Mp9@1343_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1342 N_OUT9_Mp9@1342_d N_OUT8_Mp9@1342_g N_VDD_Mp9@1342_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1341 N_OUT9_Mn9@1341_d N_OUT8_Mn9@1341_g N_VSS_Mn9@1341_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1340 N_OUT9_Mn9@1340_d N_OUT8_Mn9@1340_g N_VSS_Mn9@1340_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1341 N_OUT9_Mp9@1341_d N_OUT8_Mp9@1341_g N_VDD_Mp9@1341_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1340 N_OUT9_Mp9@1340_d N_OUT8_Mp9@1340_g N_VDD_Mp9@1340_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1339 N_OUT9_Mn9@1339_d N_OUT8_Mn9@1339_g N_VSS_Mn9@1339_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1338 N_OUT9_Mn9@1338_d N_OUT8_Mn9@1338_g N_VSS_Mn9@1338_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1339 N_OUT9_Mp9@1339_d N_OUT8_Mp9@1339_g N_VDD_Mp9@1339_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1338 N_OUT9_Mp9@1338_d N_OUT8_Mp9@1338_g N_VDD_Mp9@1338_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1337 N_OUT9_Mn9@1337_d N_OUT8_Mn9@1337_g N_VSS_Mn9@1337_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1336 N_OUT9_Mn9@1336_d N_OUT8_Mn9@1336_g N_VSS_Mn9@1336_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1337 N_OUT9_Mp9@1337_d N_OUT8_Mp9@1337_g N_VDD_Mp9@1337_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1336 N_OUT9_Mp9@1336_d N_OUT8_Mp9@1336_g N_VDD_Mp9@1336_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1335 N_OUT9_Mn9@1335_d N_OUT8_Mn9@1335_g N_VSS_Mn9@1335_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1334 N_OUT9_Mn9@1334_d N_OUT8_Mn9@1334_g N_VSS_Mn9@1334_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1335 N_OUT9_Mp9@1335_d N_OUT8_Mp9@1335_g N_VDD_Mp9@1335_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1334 N_OUT9_Mp9@1334_d N_OUT8_Mp9@1334_g N_VDD_Mp9@1334_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1333 N_OUT9_Mn9@1333_d N_OUT8_Mn9@1333_g N_VSS_Mn9@1333_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1332 N_OUT9_Mn9@1332_d N_OUT8_Mn9@1332_g N_VSS_Mn9@1332_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1333 N_OUT9_Mp9@1333_d N_OUT8_Mp9@1333_g N_VDD_Mp9@1333_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1332 N_OUT9_Mp9@1332_d N_OUT8_Mp9@1332_g N_VDD_Mp9@1332_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1331 N_OUT9_Mn9@1331_d N_OUT8_Mn9@1331_g N_VSS_Mn9@1331_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1330 N_OUT9_Mn9@1330_d N_OUT8_Mn9@1330_g N_VSS_Mn9@1330_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1331 N_OUT9_Mp9@1331_d N_OUT8_Mp9@1331_g N_VDD_Mp9@1331_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1330 N_OUT9_Mp9@1330_d N_OUT8_Mp9@1330_g N_VDD_Mp9@1330_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1329 N_OUT9_Mn9@1329_d N_OUT8_Mn9@1329_g N_VSS_Mn9@1329_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1328 N_OUT9_Mn9@1328_d N_OUT8_Mn9@1328_g N_VSS_Mn9@1328_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1329 N_OUT9_Mp9@1329_d N_OUT8_Mp9@1329_g N_VDD_Mp9@1329_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1328 N_OUT9_Mp9@1328_d N_OUT8_Mp9@1328_g N_VDD_Mp9@1328_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1327 N_OUT9_Mn9@1327_d N_OUT8_Mn9@1327_g N_VSS_Mn9@1327_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1326 N_OUT9_Mn9@1326_d N_OUT8_Mn9@1326_g N_VSS_Mn9@1326_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1327 N_OUT9_Mp9@1327_d N_OUT8_Mp9@1327_g N_VDD_Mp9@1327_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1326 N_OUT9_Mp9@1326_d N_OUT8_Mp9@1326_g N_VDD_Mp9@1326_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1325 N_OUT9_Mn9@1325_d N_OUT8_Mn9@1325_g N_VSS_Mn9@1325_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1324 N_OUT9_Mn9@1324_d N_OUT8_Mn9@1324_g N_VSS_Mn9@1324_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1325 N_OUT9_Mp9@1325_d N_OUT8_Mp9@1325_g N_VDD_Mp9@1325_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1324 N_OUT9_Mp9@1324_d N_OUT8_Mp9@1324_g N_VDD_Mp9@1324_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1323 N_OUT9_Mn9@1323_d N_OUT8_Mn9@1323_g N_VSS_Mn9@1323_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1322 N_OUT9_Mn9@1322_d N_OUT8_Mn9@1322_g N_VSS_Mn9@1322_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1323 N_OUT9_Mp9@1323_d N_OUT8_Mp9@1323_g N_VDD_Mp9@1323_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1322 N_OUT9_Mp9@1322_d N_OUT8_Mp9@1322_g N_VDD_Mp9@1322_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1321 N_OUT9_Mn9@1321_d N_OUT8_Mn9@1321_g N_VSS_Mn9@1321_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1320 N_OUT9_Mn9@1320_d N_OUT8_Mn9@1320_g N_VSS_Mn9@1320_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1321 N_OUT9_Mp9@1321_d N_OUT8_Mp9@1321_g N_VDD_Mp9@1321_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1320 N_OUT9_Mp9@1320_d N_OUT8_Mp9@1320_g N_VDD_Mp9@1320_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1319 N_OUT9_Mn9@1319_d N_OUT8_Mn9@1319_g N_VSS_Mn9@1319_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1318 N_OUT9_Mn9@1318_d N_OUT8_Mn9@1318_g N_VSS_Mn9@1318_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1319 N_OUT9_Mp9@1319_d N_OUT8_Mp9@1319_g N_VDD_Mp9@1319_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1318 N_OUT9_Mp9@1318_d N_OUT8_Mp9@1318_g N_VDD_Mp9@1318_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1317 N_OUT9_Mn9@1317_d N_OUT8_Mn9@1317_g N_VSS_Mn9@1317_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1316 N_OUT9_Mn9@1316_d N_OUT8_Mn9@1316_g N_VSS_Mn9@1316_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1317 N_OUT9_Mp9@1317_d N_OUT8_Mp9@1317_g N_VDD_Mp9@1317_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1316 N_OUT9_Mp9@1316_d N_OUT8_Mp9@1316_g N_VDD_Mp9@1316_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1315 N_OUT9_Mn9@1315_d N_OUT8_Mn9@1315_g N_VSS_Mn9@1315_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1314 N_OUT9_Mn9@1314_d N_OUT8_Mn9@1314_g N_VSS_Mn9@1314_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1315 N_OUT9_Mp9@1315_d N_OUT8_Mp9@1315_g N_VDD_Mp9@1315_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1314 N_OUT9_Mp9@1314_d N_OUT8_Mp9@1314_g N_VDD_Mp9@1314_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1313 N_OUT9_Mn9@1313_d N_OUT8_Mn9@1313_g N_VSS_Mn9@1313_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1312 N_OUT9_Mn9@1312_d N_OUT8_Mn9@1312_g N_VSS_Mn9@1312_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1313 N_OUT9_Mp9@1313_d N_OUT8_Mp9@1313_g N_VDD_Mp9@1313_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1312 N_OUT9_Mp9@1312_d N_OUT8_Mp9@1312_g N_VDD_Mp9@1312_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1311 N_OUT9_Mn9@1311_d N_OUT8_Mn9@1311_g N_VSS_Mn9@1311_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1310 N_OUT9_Mn9@1310_d N_OUT8_Mn9@1310_g N_VSS_Mn9@1310_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1311 N_OUT9_Mp9@1311_d N_OUT8_Mp9@1311_g N_VDD_Mp9@1311_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1310 N_OUT9_Mp9@1310_d N_OUT8_Mp9@1310_g N_VDD_Mp9@1310_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1309 N_OUT9_Mn9@1309_d N_OUT8_Mn9@1309_g N_VSS_Mn9@1309_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1308 N_OUT9_Mn9@1308_d N_OUT8_Mn9@1308_g N_VSS_Mn9@1308_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1309 N_OUT9_Mp9@1309_d N_OUT8_Mp9@1309_g N_VDD_Mp9@1309_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1308 N_OUT9_Mp9@1308_d N_OUT8_Mp9@1308_g N_VDD_Mp9@1308_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1307 N_OUT9_Mn9@1307_d N_OUT8_Mn9@1307_g N_VSS_Mn9@1307_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1306 N_OUT9_Mn9@1306_d N_OUT8_Mn9@1306_g N_VSS_Mn9@1306_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1307 N_OUT9_Mp9@1307_d N_OUT8_Mp9@1307_g N_VDD_Mp9@1307_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1306 N_OUT9_Mp9@1306_d N_OUT8_Mp9@1306_g N_VDD_Mp9@1306_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1305 N_OUT9_Mn9@1305_d N_OUT8_Mn9@1305_g N_VSS_Mn9@1305_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1304 N_OUT9_Mn9@1304_d N_OUT8_Mn9@1304_g N_VSS_Mn9@1304_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1305 N_OUT9_Mp9@1305_d N_OUT8_Mp9@1305_g N_VDD_Mp9@1305_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1304 N_OUT9_Mp9@1304_d N_OUT8_Mp9@1304_g N_VDD_Mp9@1304_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1303 N_OUT9_Mn9@1303_d N_OUT8_Mn9@1303_g N_VSS_Mn9@1303_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1302 N_OUT9_Mn9@1302_d N_OUT8_Mn9@1302_g N_VSS_Mn9@1302_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1303 N_OUT9_Mp9@1303_d N_OUT8_Mp9@1303_g N_VDD_Mp9@1303_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1302 N_OUT9_Mp9@1302_d N_OUT8_Mp9@1302_g N_VDD_Mp9@1302_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1301 N_OUT9_Mn9@1301_d N_OUT8_Mn9@1301_g N_VSS_Mn9@1301_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1300 N_OUT9_Mn9@1300_d N_OUT8_Mn9@1300_g N_VSS_Mn9@1300_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1301 N_OUT9_Mp9@1301_d N_OUT8_Mp9@1301_g N_VDD_Mp9@1301_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1300 N_OUT9_Mp9@1300_d N_OUT8_Mp9@1300_g N_VDD_Mp9@1300_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1299 N_OUT9_Mn9@1299_d N_OUT8_Mn9@1299_g N_VSS_Mn9@1299_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1298 N_OUT9_Mn9@1298_d N_OUT8_Mn9@1298_g N_VSS_Mn9@1298_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1299 N_OUT9_Mp9@1299_d N_OUT8_Mp9@1299_g N_VDD_Mp9@1299_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1298 N_OUT9_Mp9@1298_d N_OUT8_Mp9@1298_g N_VDD_Mp9@1298_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1297 N_OUT9_Mn9@1297_d N_OUT8_Mn9@1297_g N_VSS_Mn9@1297_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1296 N_OUT9_Mn9@1296_d N_OUT8_Mn9@1296_g N_VSS_Mn9@1296_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1297 N_OUT9_Mp9@1297_d N_OUT8_Mp9@1297_g N_VDD_Mp9@1297_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1296 N_OUT9_Mp9@1296_d N_OUT8_Mp9@1296_g N_VDD_Mp9@1296_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1295 N_OUT9_Mn9@1295_d N_OUT8_Mn9@1295_g N_VSS_Mn9@1295_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1294 N_OUT9_Mn9@1294_d N_OUT8_Mn9@1294_g N_VSS_Mn9@1294_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1295 N_OUT9_Mp9@1295_d N_OUT8_Mp9@1295_g N_VDD_Mp9@1295_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1294 N_OUT9_Mp9@1294_d N_OUT8_Mp9@1294_g N_VDD_Mp9@1294_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1293 N_OUT9_Mn9@1293_d N_OUT8_Mn9@1293_g N_VSS_Mn9@1293_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1292 N_OUT9_Mn9@1292_d N_OUT8_Mn9@1292_g N_VSS_Mn9@1292_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1293 N_OUT9_Mp9@1293_d N_OUT8_Mp9@1293_g N_VDD_Mp9@1293_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1292 N_OUT9_Mp9@1292_d N_OUT8_Mp9@1292_g N_VDD_Mp9@1292_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1291 N_OUT9_Mn9@1291_d N_OUT8_Mn9@1291_g N_VSS_Mn9@1291_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1290 N_OUT9_Mn9@1290_d N_OUT8_Mn9@1290_g N_VSS_Mn9@1290_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1291 N_OUT9_Mp9@1291_d N_OUT8_Mp9@1291_g N_VDD_Mp9@1291_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1290 N_OUT9_Mp9@1290_d N_OUT8_Mp9@1290_g N_VDD_Mp9@1290_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1289 N_OUT9_Mn9@1289_d N_OUT8_Mn9@1289_g N_VSS_Mn9@1289_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1288 N_OUT9_Mn9@1288_d N_OUT8_Mn9@1288_g N_VSS_Mn9@1288_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1289 N_OUT9_Mp9@1289_d N_OUT8_Mp9@1289_g N_VDD_Mp9@1289_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1288 N_OUT9_Mp9@1288_d N_OUT8_Mp9@1288_g N_VDD_Mp9@1288_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1287 N_OUT9_Mn9@1287_d N_OUT8_Mn9@1287_g N_VSS_Mn9@1287_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1286 N_OUT9_Mn9@1286_d N_OUT8_Mn9@1286_g N_VSS_Mn9@1286_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1287 N_OUT9_Mp9@1287_d N_OUT8_Mp9@1287_g N_VDD_Mp9@1287_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1286 N_OUT9_Mp9@1286_d N_OUT8_Mp9@1286_g N_VDD_Mp9@1286_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1285 N_OUT9_Mn9@1285_d N_OUT8_Mn9@1285_g N_VSS_Mn9@1285_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1284 N_OUT9_Mn9@1284_d N_OUT8_Mn9@1284_g N_VSS_Mn9@1284_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1285 N_OUT9_Mp9@1285_d N_OUT8_Mp9@1285_g N_VDD_Mp9@1285_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1284 N_OUT9_Mp9@1284_d N_OUT8_Mp9@1284_g N_VDD_Mp9@1284_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1283 N_OUT9_Mn9@1283_d N_OUT8_Mn9@1283_g N_VSS_Mn9@1283_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1282 N_OUT9_Mn9@1282_d N_OUT8_Mn9@1282_g N_VSS_Mn9@1282_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1283 N_OUT9_Mp9@1283_d N_OUT8_Mp9@1283_g N_VDD_Mp9@1283_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1282 N_OUT9_Mp9@1282_d N_OUT8_Mp9@1282_g N_VDD_Mp9@1282_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1281 N_OUT9_Mn9@1281_d N_OUT8_Mn9@1281_g N_VSS_Mn9@1281_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1280 N_OUT9_Mn9@1280_d N_OUT8_Mn9@1280_g N_VSS_Mn9@1280_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1281 N_OUT9_Mp9@1281_d N_OUT8_Mp9@1281_g N_VDD_Mp9@1281_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1280 N_OUT9_Mp9@1280_d N_OUT8_Mp9@1280_g N_VDD_Mp9@1280_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1279 N_OUT9_Mn9@1279_d N_OUT8_Mn9@1279_g N_VSS_Mn9@1279_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1278 N_OUT9_Mn9@1278_d N_OUT8_Mn9@1278_g N_VSS_Mn9@1278_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1279 N_OUT9_Mp9@1279_d N_OUT8_Mp9@1279_g N_VDD_Mp9@1279_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1278 N_OUT9_Mp9@1278_d N_OUT8_Mp9@1278_g N_VDD_Mp9@1278_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1277 N_OUT9_Mn9@1277_d N_OUT8_Mn9@1277_g N_VSS_Mn9@1277_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1276 N_OUT9_Mn9@1276_d N_OUT8_Mn9@1276_g N_VSS_Mn9@1276_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1277 N_OUT9_Mp9@1277_d N_OUT8_Mp9@1277_g N_VDD_Mp9@1277_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1276 N_OUT9_Mp9@1276_d N_OUT8_Mp9@1276_g N_VDD_Mp9@1276_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1275 N_OUT9_Mn9@1275_d N_OUT8_Mn9@1275_g N_VSS_Mn9@1275_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1274 N_OUT9_Mn9@1274_d N_OUT8_Mn9@1274_g N_VSS_Mn9@1274_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1275 N_OUT9_Mp9@1275_d N_OUT8_Mp9@1275_g N_VDD_Mp9@1275_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1274 N_OUT9_Mp9@1274_d N_OUT8_Mp9@1274_g N_VDD_Mp9@1274_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1273 N_OUT9_Mn9@1273_d N_OUT8_Mn9@1273_g N_VSS_Mn9@1273_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1272 N_OUT9_Mn9@1272_d N_OUT8_Mn9@1272_g N_VSS_Mn9@1272_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1273 N_OUT9_Mp9@1273_d N_OUT8_Mp9@1273_g N_VDD_Mp9@1273_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1272 N_OUT9_Mp9@1272_d N_OUT8_Mp9@1272_g N_VDD_Mp9@1272_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1271 N_OUT9_Mn9@1271_d N_OUT8_Mn9@1271_g N_VSS_Mn9@1271_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1270 N_OUT9_Mn9@1270_d N_OUT8_Mn9@1270_g N_VSS_Mn9@1270_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1271 N_OUT9_Mp9@1271_d N_OUT8_Mp9@1271_g N_VDD_Mp9@1271_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1270 N_OUT9_Mp9@1270_d N_OUT8_Mp9@1270_g N_VDD_Mp9@1270_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1269 N_OUT9_Mn9@1269_d N_OUT8_Mn9@1269_g N_VSS_Mn9@1269_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1268 N_OUT9_Mn9@1268_d N_OUT8_Mn9@1268_g N_VSS_Mn9@1268_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1269 N_OUT9_Mp9@1269_d N_OUT8_Mp9@1269_g N_VDD_Mp9@1269_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1268 N_OUT9_Mp9@1268_d N_OUT8_Mp9@1268_g N_VDD_Mp9@1268_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1267 N_OUT9_Mn9@1267_d N_OUT8_Mn9@1267_g N_VSS_Mn9@1267_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1266 N_OUT9_Mn9@1266_d N_OUT8_Mn9@1266_g N_VSS_Mn9@1266_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1267 N_OUT9_Mp9@1267_d N_OUT8_Mp9@1267_g N_VDD_Mp9@1267_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1266 N_OUT9_Mp9@1266_d N_OUT8_Mp9@1266_g N_VDD_Mp9@1266_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1265 N_OUT9_Mn9@1265_d N_OUT8_Mn9@1265_g N_VSS_Mn9@1265_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1264 N_OUT9_Mn9@1264_d N_OUT8_Mn9@1264_g N_VSS_Mn9@1264_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1265 N_OUT9_Mp9@1265_d N_OUT8_Mp9@1265_g N_VDD_Mp9@1265_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1264 N_OUT9_Mp9@1264_d N_OUT8_Mp9@1264_g N_VDD_Mp9@1264_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1263 N_OUT9_Mn9@1263_d N_OUT8_Mn9@1263_g N_VSS_Mn9@1263_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1262 N_OUT9_Mn9@1262_d N_OUT8_Mn9@1262_g N_VSS_Mn9@1262_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1263 N_OUT9_Mp9@1263_d N_OUT8_Mp9@1263_g N_VDD_Mp9@1263_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1262 N_OUT9_Mp9@1262_d N_OUT8_Mp9@1262_g N_VDD_Mp9@1262_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1261 N_OUT9_Mn9@1261_d N_OUT8_Mn9@1261_g N_VSS_Mn9@1261_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1260 N_OUT9_Mn9@1260_d N_OUT8_Mn9@1260_g N_VSS_Mn9@1260_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1261 N_OUT9_Mp9@1261_d N_OUT8_Mp9@1261_g N_VDD_Mp9@1261_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1260 N_OUT9_Mp9@1260_d N_OUT8_Mp9@1260_g N_VDD_Mp9@1260_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1259 N_OUT9_Mn9@1259_d N_OUT8_Mn9@1259_g N_VSS_Mn9@1259_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1258 N_OUT9_Mn9@1258_d N_OUT8_Mn9@1258_g N_VSS_Mn9@1258_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1259 N_OUT9_Mp9@1259_d N_OUT8_Mp9@1259_g N_VDD_Mp9@1259_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1258 N_OUT9_Mp9@1258_d N_OUT8_Mp9@1258_g N_VDD_Mp9@1258_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1257 N_OUT9_Mn9@1257_d N_OUT8_Mn9@1257_g N_VSS_Mn9@1257_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1256 N_OUT9_Mn9@1256_d N_OUT8_Mn9@1256_g N_VSS_Mn9@1256_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1257 N_OUT9_Mp9@1257_d N_OUT8_Mp9@1257_g N_VDD_Mp9@1257_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1256 N_OUT9_Mp9@1256_d N_OUT8_Mp9@1256_g N_VDD_Mp9@1256_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1255 N_OUT9_Mn9@1255_d N_OUT8_Mn9@1255_g N_VSS_Mn9@1255_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1254 N_OUT9_Mn9@1254_d N_OUT8_Mn9@1254_g N_VSS_Mn9@1254_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1255 N_OUT9_Mp9@1255_d N_OUT8_Mp9@1255_g N_VDD_Mp9@1255_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1254 N_OUT9_Mp9@1254_d N_OUT8_Mp9@1254_g N_VDD_Mp9@1254_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1253 N_OUT9_Mn9@1253_d N_OUT8_Mn9@1253_g N_VSS_Mn9@1253_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1252 N_OUT9_Mn9@1252_d N_OUT8_Mn9@1252_g N_VSS_Mn9@1252_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1253 N_OUT9_Mp9@1253_d N_OUT8_Mp9@1253_g N_VDD_Mp9@1253_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1252 N_OUT9_Mp9@1252_d N_OUT8_Mp9@1252_g N_VDD_Mp9@1252_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1251 N_OUT9_Mn9@1251_d N_OUT8_Mn9@1251_g N_VSS_Mn9@1251_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1250 N_OUT9_Mn9@1250_d N_OUT8_Mn9@1250_g N_VSS_Mn9@1250_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1251 N_OUT9_Mp9@1251_d N_OUT8_Mp9@1251_g N_VDD_Mp9@1251_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1250 N_OUT9_Mp9@1250_d N_OUT8_Mp9@1250_g N_VDD_Mp9@1250_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1249 N_OUT9_Mn9@1249_d N_OUT8_Mn9@1249_g N_VSS_Mn9@1249_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1248 N_OUT9_Mn9@1248_d N_OUT8_Mn9@1248_g N_VSS_Mn9@1248_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1249 N_OUT9_Mp9@1249_d N_OUT8_Mp9@1249_g N_VDD_Mp9@1249_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1248 N_OUT9_Mp9@1248_d N_OUT8_Mp9@1248_g N_VDD_Mp9@1248_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1247 N_OUT9_Mn9@1247_d N_OUT8_Mn9@1247_g N_VSS_Mn9@1247_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1246 N_OUT9_Mn9@1246_d N_OUT8_Mn9@1246_g N_VSS_Mn9@1246_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1247 N_OUT9_Mp9@1247_d N_OUT8_Mp9@1247_g N_VDD_Mp9@1247_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1246 N_OUT9_Mp9@1246_d N_OUT8_Mp9@1246_g N_VDD_Mp9@1246_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1245 N_OUT9_Mn9@1245_d N_OUT8_Mn9@1245_g N_VSS_Mn9@1245_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1244 N_OUT9_Mn9@1244_d N_OUT8_Mn9@1244_g N_VSS_Mn9@1244_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1245 N_OUT9_Mp9@1245_d N_OUT8_Mp9@1245_g N_VDD_Mp9@1245_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1244 N_OUT9_Mp9@1244_d N_OUT8_Mp9@1244_g N_VDD_Mp9@1244_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1243 N_OUT9_Mn9@1243_d N_OUT8_Mn9@1243_g N_VSS_Mn9@1243_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1242 N_OUT9_Mn9@1242_d N_OUT8_Mn9@1242_g N_VSS_Mn9@1242_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1243 N_OUT9_Mp9@1243_d N_OUT8_Mp9@1243_g N_VDD_Mp9@1243_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1242 N_OUT9_Mp9@1242_d N_OUT8_Mp9@1242_g N_VDD_Mp9@1242_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1241 N_OUT9_Mn9@1241_d N_OUT8_Mn9@1241_g N_VSS_Mn9@1241_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1240 N_OUT9_Mn9@1240_d N_OUT8_Mn9@1240_g N_VSS_Mn9@1240_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1241 N_OUT9_Mp9@1241_d N_OUT8_Mp9@1241_g N_VDD_Mp9@1241_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1240 N_OUT9_Mp9@1240_d N_OUT8_Mp9@1240_g N_VDD_Mp9@1240_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1239 N_OUT9_Mn9@1239_d N_OUT8_Mn9@1239_g N_VSS_Mn9@1239_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1238 N_OUT9_Mn9@1238_d N_OUT8_Mn9@1238_g N_VSS_Mn9@1238_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1239 N_OUT9_Mp9@1239_d N_OUT8_Mp9@1239_g N_VDD_Mp9@1239_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1238 N_OUT9_Mp9@1238_d N_OUT8_Mp9@1238_g N_VDD_Mp9@1238_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1237 N_OUT9_Mn9@1237_d N_OUT8_Mn9@1237_g N_VSS_Mn9@1237_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1236 N_OUT9_Mn9@1236_d N_OUT8_Mn9@1236_g N_VSS_Mn9@1236_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1237 N_OUT9_Mp9@1237_d N_OUT8_Mp9@1237_g N_VDD_Mp9@1237_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1236 N_OUT9_Mp9@1236_d N_OUT8_Mp9@1236_g N_VDD_Mp9@1236_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1235 N_OUT9_Mn9@1235_d N_OUT8_Mn9@1235_g N_VSS_Mn9@1235_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1234 N_OUT9_Mn9@1234_d N_OUT8_Mn9@1234_g N_VSS_Mn9@1234_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1235 N_OUT9_Mp9@1235_d N_OUT8_Mp9@1235_g N_VDD_Mp9@1235_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1234 N_OUT9_Mp9@1234_d N_OUT8_Mp9@1234_g N_VDD_Mp9@1234_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1233 N_OUT9_Mn9@1233_d N_OUT8_Mn9@1233_g N_VSS_Mn9@1233_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1232 N_OUT9_Mn9@1232_d N_OUT8_Mn9@1232_g N_VSS_Mn9@1232_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1233 N_OUT9_Mp9@1233_d N_OUT8_Mp9@1233_g N_VDD_Mp9@1233_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1232 N_OUT9_Mp9@1232_d N_OUT8_Mp9@1232_g N_VDD_Mp9@1232_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1231 N_OUT9_Mn9@1231_d N_OUT8_Mn9@1231_g N_VSS_Mn9@1231_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1230 N_OUT9_Mn9@1230_d N_OUT8_Mn9@1230_g N_VSS_Mn9@1230_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1231 N_OUT9_Mp9@1231_d N_OUT8_Mp9@1231_g N_VDD_Mp9@1231_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1230 N_OUT9_Mp9@1230_d N_OUT8_Mp9@1230_g N_VDD_Mp9@1230_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1229 N_OUT9_Mn9@1229_d N_OUT8_Mn9@1229_g N_VSS_Mn9@1229_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1228 N_OUT9_Mn9@1228_d N_OUT8_Mn9@1228_g N_VSS_Mn9@1228_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1229 N_OUT9_Mp9@1229_d N_OUT8_Mp9@1229_g N_VDD_Mp9@1229_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1228 N_OUT9_Mp9@1228_d N_OUT8_Mp9@1228_g N_VDD_Mp9@1228_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1227 N_OUT9_Mn9@1227_d N_OUT8_Mn9@1227_g N_VSS_Mn9@1227_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1226 N_OUT9_Mn9@1226_d N_OUT8_Mn9@1226_g N_VSS_Mn9@1226_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1227 N_OUT9_Mp9@1227_d N_OUT8_Mp9@1227_g N_VDD_Mp9@1227_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1226 N_OUT9_Mp9@1226_d N_OUT8_Mp9@1226_g N_VDD_Mp9@1226_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1225 N_OUT9_Mn9@1225_d N_OUT8_Mn9@1225_g N_VSS_Mn9@1225_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1224 N_OUT9_Mn9@1224_d N_OUT8_Mn9@1224_g N_VSS_Mn9@1224_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1225 N_OUT9_Mp9@1225_d N_OUT8_Mp9@1225_g N_VDD_Mp9@1225_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1224 N_OUT9_Mp9@1224_d N_OUT8_Mp9@1224_g N_VDD_Mp9@1224_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1223 N_OUT9_Mn9@1223_d N_OUT8_Mn9@1223_g N_VSS_Mn9@1223_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1222 N_OUT9_Mn9@1222_d N_OUT8_Mn9@1222_g N_VSS_Mn9@1222_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1223 N_OUT9_Mp9@1223_d N_OUT8_Mp9@1223_g N_VDD_Mp9@1223_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1222 N_OUT9_Mp9@1222_d N_OUT8_Mp9@1222_g N_VDD_Mp9@1222_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1221 N_OUT9_Mn9@1221_d N_OUT8_Mn9@1221_g N_VSS_Mn9@1221_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1220 N_OUT9_Mn9@1220_d N_OUT8_Mn9@1220_g N_VSS_Mn9@1220_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1221 N_OUT9_Mp9@1221_d N_OUT8_Mp9@1221_g N_VDD_Mp9@1221_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1220 N_OUT9_Mp9@1220_d N_OUT8_Mp9@1220_g N_VDD_Mp9@1220_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1219 N_OUT9_Mn9@1219_d N_OUT8_Mn9@1219_g N_VSS_Mn9@1219_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1218 N_OUT9_Mn9@1218_d N_OUT8_Mn9@1218_g N_VSS_Mn9@1218_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1219 N_OUT9_Mp9@1219_d N_OUT8_Mp9@1219_g N_VDD_Mp9@1219_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1218 N_OUT9_Mp9@1218_d N_OUT8_Mp9@1218_g N_VDD_Mp9@1218_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1217 N_OUT9_Mn9@1217_d N_OUT8_Mn9@1217_g N_VSS_Mn9@1217_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1216 N_OUT9_Mn9@1216_d N_OUT8_Mn9@1216_g N_VSS_Mn9@1216_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1217 N_OUT9_Mp9@1217_d N_OUT8_Mp9@1217_g N_VDD_Mp9@1217_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1216 N_OUT9_Mp9@1216_d N_OUT8_Mp9@1216_g N_VDD_Mp9@1216_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1215 N_OUT9_Mn9@1215_d N_OUT8_Mn9@1215_g N_VSS_Mn9@1215_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1214 N_OUT9_Mn9@1214_d N_OUT8_Mn9@1214_g N_VSS_Mn9@1214_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1215 N_OUT9_Mp9@1215_d N_OUT8_Mp9@1215_g N_VDD_Mp9@1215_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1214 N_OUT9_Mp9@1214_d N_OUT8_Mp9@1214_g N_VDD_Mp9@1214_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1213 N_OUT9_Mn9@1213_d N_OUT8_Mn9@1213_g N_VSS_Mn9@1213_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1212 N_OUT9_Mn9@1212_d N_OUT8_Mn9@1212_g N_VSS_Mn9@1212_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1213 N_OUT9_Mp9@1213_d N_OUT8_Mp9@1213_g N_VDD_Mp9@1213_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1212 N_OUT9_Mp9@1212_d N_OUT8_Mp9@1212_g N_VDD_Mp9@1212_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1211 N_OUT9_Mn9@1211_d N_OUT8_Mn9@1211_g N_VSS_Mn9@1211_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1210 N_OUT9_Mn9@1210_d N_OUT8_Mn9@1210_g N_VSS_Mn9@1210_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1211 N_OUT9_Mp9@1211_d N_OUT8_Mp9@1211_g N_VDD_Mp9@1211_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1210 N_OUT9_Mp9@1210_d N_OUT8_Mp9@1210_g N_VDD_Mp9@1210_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1209 N_OUT9_Mn9@1209_d N_OUT8_Mn9@1209_g N_VSS_Mn9@1209_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1208 N_OUT9_Mn9@1208_d N_OUT8_Mn9@1208_g N_VSS_Mn9@1208_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1209 N_OUT9_Mp9@1209_d N_OUT8_Mp9@1209_g N_VDD_Mp9@1209_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1208 N_OUT9_Mp9@1208_d N_OUT8_Mp9@1208_g N_VDD_Mp9@1208_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1207 N_OUT9_Mn9@1207_d N_OUT8_Mn9@1207_g N_VSS_Mn9@1207_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1206 N_OUT9_Mn9@1206_d N_OUT8_Mn9@1206_g N_VSS_Mn9@1206_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1207 N_OUT9_Mp9@1207_d N_OUT8_Mp9@1207_g N_VDD_Mp9@1207_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1206 N_OUT9_Mp9@1206_d N_OUT8_Mp9@1206_g N_VDD_Mp9@1206_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1205 N_OUT9_Mn9@1205_d N_OUT8_Mn9@1205_g N_VSS_Mn9@1205_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1204 N_OUT9_Mn9@1204_d N_OUT8_Mn9@1204_g N_VSS_Mn9@1204_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1205 N_OUT9_Mp9@1205_d N_OUT8_Mp9@1205_g N_VDD_Mp9@1205_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1204 N_OUT9_Mp9@1204_d N_OUT8_Mp9@1204_g N_VDD_Mp9@1204_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1203 N_OUT9_Mn9@1203_d N_OUT8_Mn9@1203_g N_VSS_Mn9@1203_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1202 N_OUT9_Mn9@1202_d N_OUT8_Mn9@1202_g N_VSS_Mn9@1202_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1203 N_OUT9_Mp9@1203_d N_OUT8_Mp9@1203_g N_VDD_Mp9@1203_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1202 N_OUT9_Mp9@1202_d N_OUT8_Mp9@1202_g N_VDD_Mp9@1202_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1201 N_OUT9_Mn9@1201_d N_OUT8_Mn9@1201_g N_VSS_Mn9@1201_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1200 N_OUT9_Mn9@1200_d N_OUT8_Mn9@1200_g N_VSS_Mn9@1200_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1201 N_OUT9_Mp9@1201_d N_OUT8_Mp9@1201_g N_VDD_Mp9@1201_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1200 N_OUT9_Mp9@1200_d N_OUT8_Mp9@1200_g N_VDD_Mp9@1200_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1199 N_OUT9_Mn9@1199_d N_OUT8_Mn9@1199_g N_VSS_Mn9@1199_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1198 N_OUT9_Mn9@1198_d N_OUT8_Mn9@1198_g N_VSS_Mn9@1198_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1199 N_OUT9_Mp9@1199_d N_OUT8_Mp9@1199_g N_VDD_Mp9@1199_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1198 N_OUT9_Mp9@1198_d N_OUT8_Mp9@1198_g N_VDD_Mp9@1198_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1197 N_OUT9_Mn9@1197_d N_OUT8_Mn9@1197_g N_VSS_Mn9@1197_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1196 N_OUT9_Mn9@1196_d N_OUT8_Mn9@1196_g N_VSS_Mn9@1196_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1197 N_OUT9_Mp9@1197_d N_OUT8_Mp9@1197_g N_VDD_Mp9@1197_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1196 N_OUT9_Mp9@1196_d N_OUT8_Mp9@1196_g N_VDD_Mp9@1196_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1195 N_OUT9_Mn9@1195_d N_OUT8_Mn9@1195_g N_VSS_Mn9@1195_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1194 N_OUT9_Mn9@1194_d N_OUT8_Mn9@1194_g N_VSS_Mn9@1194_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1195 N_OUT9_Mp9@1195_d N_OUT8_Mp9@1195_g N_VDD_Mp9@1195_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1194 N_OUT9_Mp9@1194_d N_OUT8_Mp9@1194_g N_VDD_Mp9@1194_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1193 N_OUT9_Mn9@1193_d N_OUT8_Mn9@1193_g N_VSS_Mn9@1193_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1192 N_OUT9_Mn9@1192_d N_OUT8_Mn9@1192_g N_VSS_Mn9@1192_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1193 N_OUT9_Mp9@1193_d N_OUT8_Mp9@1193_g N_VDD_Mp9@1193_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1192 N_OUT9_Mp9@1192_d N_OUT8_Mp9@1192_g N_VDD_Mp9@1192_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1191 N_OUT9_Mn9@1191_d N_OUT8_Mn9@1191_g N_VSS_Mn9@1191_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1190 N_OUT9_Mn9@1190_d N_OUT8_Mn9@1190_g N_VSS_Mn9@1190_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1191 N_OUT9_Mp9@1191_d N_OUT8_Mp9@1191_g N_VDD_Mp9@1191_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1190 N_OUT9_Mp9@1190_d N_OUT8_Mp9@1190_g N_VDD_Mp9@1190_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1189 N_OUT9_Mn9@1189_d N_OUT8_Mn9@1189_g N_VSS_Mn9@1189_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1188 N_OUT9_Mn9@1188_d N_OUT8_Mn9@1188_g N_VSS_Mn9@1188_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1189 N_OUT9_Mp9@1189_d N_OUT8_Mp9@1189_g N_VDD_Mp9@1189_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1188 N_OUT9_Mp9@1188_d N_OUT8_Mp9@1188_g N_VDD_Mp9@1188_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1187 N_OUT9_Mn9@1187_d N_OUT8_Mn9@1187_g N_VSS_Mn9@1187_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1186 N_OUT9_Mn9@1186_d N_OUT8_Mn9@1186_g N_VSS_Mn9@1186_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1187 N_OUT9_Mp9@1187_d N_OUT8_Mp9@1187_g N_VDD_Mp9@1187_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1186 N_OUT9_Mp9@1186_d N_OUT8_Mp9@1186_g N_VDD_Mp9@1186_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1185 N_OUT9_Mn9@1185_d N_OUT8_Mn9@1185_g N_VSS_Mn9@1185_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1184 N_OUT9_Mn9@1184_d N_OUT8_Mn9@1184_g N_VSS_Mn9@1184_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1185 N_OUT9_Mp9@1185_d N_OUT8_Mp9@1185_g N_VDD_Mp9@1185_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1184 N_OUT9_Mp9@1184_d N_OUT8_Mp9@1184_g N_VDD_Mp9@1184_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1183 N_OUT9_Mn9@1183_d N_OUT8_Mn9@1183_g N_VSS_Mn9@1183_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1182 N_OUT9_Mn9@1182_d N_OUT8_Mn9@1182_g N_VSS_Mn9@1182_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1183 N_OUT9_Mp9@1183_d N_OUT8_Mp9@1183_g N_VDD_Mp9@1183_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1182 N_OUT9_Mp9@1182_d N_OUT8_Mp9@1182_g N_VDD_Mp9@1182_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1181 N_OUT9_Mn9@1181_d N_OUT8_Mn9@1181_g N_VSS_Mn9@1181_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1180 N_OUT9_Mn9@1180_d N_OUT8_Mn9@1180_g N_VSS_Mn9@1180_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1181 N_OUT9_Mp9@1181_d N_OUT8_Mp9@1181_g N_VDD_Mp9@1181_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1180 N_OUT9_Mp9@1180_d N_OUT8_Mp9@1180_g N_VDD_Mp9@1180_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1179 N_OUT9_Mn9@1179_d N_OUT8_Mn9@1179_g N_VSS_Mn9@1179_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1178 N_OUT9_Mn9@1178_d N_OUT8_Mn9@1178_g N_VSS_Mn9@1178_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1179 N_OUT9_Mp9@1179_d N_OUT8_Mp9@1179_g N_VDD_Mp9@1179_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1178 N_OUT9_Mp9@1178_d N_OUT8_Mp9@1178_g N_VDD_Mp9@1178_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1177 N_OUT9_Mn9@1177_d N_OUT8_Mn9@1177_g N_VSS_Mn9@1177_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1176 N_OUT9_Mn9@1176_d N_OUT8_Mn9@1176_g N_VSS_Mn9@1176_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1177 N_OUT9_Mp9@1177_d N_OUT8_Mp9@1177_g N_VDD_Mp9@1177_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1176 N_OUT9_Mp9@1176_d N_OUT8_Mp9@1176_g N_VDD_Mp9@1176_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1175 N_OUT9_Mn9@1175_d N_OUT8_Mn9@1175_g N_VSS_Mn9@1175_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1174 N_OUT9_Mn9@1174_d N_OUT8_Mn9@1174_g N_VSS_Mn9@1174_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1175 N_OUT9_Mp9@1175_d N_OUT8_Mp9@1175_g N_VDD_Mp9@1175_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1174 N_OUT9_Mp9@1174_d N_OUT8_Mp9@1174_g N_VDD_Mp9@1174_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1173 N_OUT9_Mn9@1173_d N_OUT8_Mn9@1173_g N_VSS_Mn9@1173_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1172 N_OUT9_Mn9@1172_d N_OUT8_Mn9@1172_g N_VSS_Mn9@1172_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1173 N_OUT9_Mp9@1173_d N_OUT8_Mp9@1173_g N_VDD_Mp9@1173_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1172 N_OUT9_Mp9@1172_d N_OUT8_Mp9@1172_g N_VDD_Mp9@1172_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1171 N_OUT9_Mn9@1171_d N_OUT8_Mn9@1171_g N_VSS_Mn9@1171_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1170 N_OUT9_Mn9@1170_d N_OUT8_Mn9@1170_g N_VSS_Mn9@1170_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1171 N_OUT9_Mp9@1171_d N_OUT8_Mp9@1171_g N_VDD_Mp9@1171_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1170 N_OUT9_Mp9@1170_d N_OUT8_Mp9@1170_g N_VDD_Mp9@1170_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1169 N_OUT9_Mn9@1169_d N_OUT8_Mn9@1169_g N_VSS_Mn9@1169_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1168 N_OUT9_Mn9@1168_d N_OUT8_Mn9@1168_g N_VSS_Mn9@1168_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1169 N_OUT9_Mp9@1169_d N_OUT8_Mp9@1169_g N_VDD_Mp9@1169_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1168 N_OUT9_Mp9@1168_d N_OUT8_Mp9@1168_g N_VDD_Mp9@1168_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1167 N_OUT9_Mn9@1167_d N_OUT8_Mn9@1167_g N_VSS_Mn9@1167_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1166 N_OUT9_Mn9@1166_d N_OUT8_Mn9@1166_g N_VSS_Mn9@1166_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1167 N_OUT9_Mp9@1167_d N_OUT8_Mp9@1167_g N_VDD_Mp9@1167_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1166 N_OUT9_Mp9@1166_d N_OUT8_Mp9@1166_g N_VDD_Mp9@1166_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1165 N_OUT9_Mn9@1165_d N_OUT8_Mn9@1165_g N_VSS_Mn9@1165_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1164 N_OUT9_Mn9@1164_d N_OUT8_Mn9@1164_g N_VSS_Mn9@1164_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1165 N_OUT9_Mp9@1165_d N_OUT8_Mp9@1165_g N_VDD_Mp9@1165_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1164 N_OUT9_Mp9@1164_d N_OUT8_Mp9@1164_g N_VDD_Mp9@1164_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1163 N_OUT9_Mn9@1163_d N_OUT8_Mn9@1163_g N_VSS_Mn9@1163_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1162 N_OUT9_Mn9@1162_d N_OUT8_Mn9@1162_g N_VSS_Mn9@1162_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1163 N_OUT9_Mp9@1163_d N_OUT8_Mp9@1163_g N_VDD_Mp9@1163_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1162 N_OUT9_Mp9@1162_d N_OUT8_Mp9@1162_g N_VDD_Mp9@1162_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1161 N_OUT9_Mn9@1161_d N_OUT8_Mn9@1161_g N_VSS_Mn9@1161_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1160 N_OUT9_Mn9@1160_d N_OUT8_Mn9@1160_g N_VSS_Mn9@1160_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1161 N_OUT9_Mp9@1161_d N_OUT8_Mp9@1161_g N_VDD_Mp9@1161_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1160 N_OUT9_Mp9@1160_d N_OUT8_Mp9@1160_g N_VDD_Mp9@1160_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1159 N_OUT9_Mn9@1159_d N_OUT8_Mn9@1159_g N_VSS_Mn9@1159_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1158 N_OUT9_Mn9@1158_d N_OUT8_Mn9@1158_g N_VSS_Mn9@1158_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1159 N_OUT9_Mp9@1159_d N_OUT8_Mp9@1159_g N_VDD_Mp9@1159_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1158 N_OUT9_Mp9@1158_d N_OUT8_Mp9@1158_g N_VDD_Mp9@1158_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1157 N_OUT9_Mn9@1157_d N_OUT8_Mn9@1157_g N_VSS_Mn9@1157_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1156 N_OUT9_Mn9@1156_d N_OUT8_Mn9@1156_g N_VSS_Mn9@1156_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1157 N_OUT9_Mp9@1157_d N_OUT8_Mp9@1157_g N_VDD_Mp9@1157_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1156 N_OUT9_Mp9@1156_d N_OUT8_Mp9@1156_g N_VDD_Mp9@1156_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1155 N_OUT9_Mn9@1155_d N_OUT8_Mn9@1155_g N_VSS_Mn9@1155_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1154 N_OUT9_Mn9@1154_d N_OUT8_Mn9@1154_g N_VSS_Mn9@1154_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1155 N_OUT9_Mp9@1155_d N_OUT8_Mp9@1155_g N_VDD_Mp9@1155_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1154 N_OUT9_Mp9@1154_d N_OUT8_Mp9@1154_g N_VDD_Mp9@1154_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1153 N_OUT9_Mn9@1153_d N_OUT8_Mn9@1153_g N_VSS_Mn9@1153_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1152 N_OUT9_Mn9@1152_d N_OUT8_Mn9@1152_g N_VSS_Mn9@1152_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1153 N_OUT9_Mp9@1153_d N_OUT8_Mp9@1153_g N_VDD_Mp9@1153_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1152 N_OUT9_Mp9@1152_d N_OUT8_Mp9@1152_g N_VDD_Mp9@1152_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1151 N_OUT9_Mn9@1151_d N_OUT8_Mn9@1151_g N_VSS_Mn9@1151_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1150 N_OUT9_Mn9@1150_d N_OUT8_Mn9@1150_g N_VSS_Mn9@1150_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1151 N_OUT9_Mp9@1151_d N_OUT8_Mp9@1151_g N_VDD_Mp9@1151_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1150 N_OUT9_Mp9@1150_d N_OUT8_Mp9@1150_g N_VDD_Mp9@1150_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1149 N_OUT9_Mn9@1149_d N_OUT8_Mn9@1149_g N_VSS_Mn9@1149_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1148 N_OUT9_Mn9@1148_d N_OUT8_Mn9@1148_g N_VSS_Mn9@1148_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1149 N_OUT9_Mp9@1149_d N_OUT8_Mp9@1149_g N_VDD_Mp9@1149_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1148 N_OUT9_Mp9@1148_d N_OUT8_Mp9@1148_g N_VDD_Mp9@1148_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1147 N_OUT9_Mn9@1147_d N_OUT8_Mn9@1147_g N_VSS_Mn9@1147_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1146 N_OUT9_Mn9@1146_d N_OUT8_Mn9@1146_g N_VSS_Mn9@1146_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1147 N_OUT9_Mp9@1147_d N_OUT8_Mp9@1147_g N_VDD_Mp9@1147_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1146 N_OUT9_Mp9@1146_d N_OUT8_Mp9@1146_g N_VDD_Mp9@1146_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1145 N_OUT9_Mn9@1145_d N_OUT8_Mn9@1145_g N_VSS_Mn9@1145_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1144 N_OUT9_Mn9@1144_d N_OUT8_Mn9@1144_g N_VSS_Mn9@1144_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1145 N_OUT9_Mp9@1145_d N_OUT8_Mp9@1145_g N_VDD_Mp9@1145_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1144 N_OUT9_Mp9@1144_d N_OUT8_Mp9@1144_g N_VDD_Mp9@1144_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1143 N_OUT9_Mn9@1143_d N_OUT8_Mn9@1143_g N_VSS_Mn9@1143_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1142 N_OUT9_Mn9@1142_d N_OUT8_Mn9@1142_g N_VSS_Mn9@1142_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1143 N_OUT9_Mp9@1143_d N_OUT8_Mp9@1143_g N_VDD_Mp9@1143_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1142 N_OUT9_Mp9@1142_d N_OUT8_Mp9@1142_g N_VDD_Mp9@1142_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1141 N_OUT9_Mn9@1141_d N_OUT8_Mn9@1141_g N_VSS_Mn9@1141_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1140 N_OUT9_Mn9@1140_d N_OUT8_Mn9@1140_g N_VSS_Mn9@1140_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1141 N_OUT9_Mp9@1141_d N_OUT8_Mp9@1141_g N_VDD_Mp9@1141_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1140 N_OUT9_Mp9@1140_d N_OUT8_Mp9@1140_g N_VDD_Mp9@1140_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1139 N_OUT9_Mn9@1139_d N_OUT8_Mn9@1139_g N_VSS_Mn9@1139_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1138 N_OUT9_Mn9@1138_d N_OUT8_Mn9@1138_g N_VSS_Mn9@1138_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1139 N_OUT9_Mp9@1139_d N_OUT8_Mp9@1139_g N_VDD_Mp9@1139_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1138 N_OUT9_Mp9@1138_d N_OUT8_Mp9@1138_g N_VDD_Mp9@1138_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1137 N_OUT9_Mn9@1137_d N_OUT8_Mn9@1137_g N_VSS_Mn9@1137_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1136 N_OUT9_Mn9@1136_d N_OUT8_Mn9@1136_g N_VSS_Mn9@1136_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1137 N_OUT9_Mp9@1137_d N_OUT8_Mp9@1137_g N_VDD_Mp9@1137_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1136 N_OUT9_Mp9@1136_d N_OUT8_Mp9@1136_g N_VDD_Mp9@1136_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1135 N_OUT9_Mn9@1135_d N_OUT8_Mn9@1135_g N_VSS_Mn9@1135_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1134 N_OUT9_Mn9@1134_d N_OUT8_Mn9@1134_g N_VSS_Mn9@1134_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1135 N_OUT9_Mp9@1135_d N_OUT8_Mp9@1135_g N_VDD_Mp9@1135_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1134 N_OUT9_Mp9@1134_d N_OUT8_Mp9@1134_g N_VDD_Mp9@1134_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1133 N_OUT9_Mn9@1133_d N_OUT8_Mn9@1133_g N_VSS_Mn9@1133_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1132 N_OUT9_Mn9@1132_d N_OUT8_Mn9@1132_g N_VSS_Mn9@1132_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1133 N_OUT9_Mp9@1133_d N_OUT8_Mp9@1133_g N_VDD_Mp9@1133_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1132 N_OUT9_Mp9@1132_d N_OUT8_Mp9@1132_g N_VDD_Mp9@1132_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1131 N_OUT9_Mn9@1131_d N_OUT8_Mn9@1131_g N_VSS_Mn9@1131_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1130 N_OUT9_Mn9@1130_d N_OUT8_Mn9@1130_g N_VSS_Mn9@1130_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1131 N_OUT9_Mp9@1131_d N_OUT8_Mp9@1131_g N_VDD_Mp9@1131_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1130 N_OUT9_Mp9@1130_d N_OUT8_Mp9@1130_g N_VDD_Mp9@1130_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1129 N_OUT9_Mn9@1129_d N_OUT8_Mn9@1129_g N_VSS_Mn9@1129_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1128 N_OUT9_Mn9@1128_d N_OUT8_Mn9@1128_g N_VSS_Mn9@1128_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1129 N_OUT9_Mp9@1129_d N_OUT8_Mp9@1129_g N_VDD_Mp9@1129_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1128 N_OUT9_Mp9@1128_d N_OUT8_Mp9@1128_g N_VDD_Mp9@1128_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1127 N_OUT9_Mn9@1127_d N_OUT8_Mn9@1127_g N_VSS_Mn9@1127_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1126 N_OUT9_Mn9@1126_d N_OUT8_Mn9@1126_g N_VSS_Mn9@1126_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1127 N_OUT9_Mp9@1127_d N_OUT8_Mp9@1127_g N_VDD_Mp9@1127_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1126 N_OUT9_Mp9@1126_d N_OUT8_Mp9@1126_g N_VDD_Mp9@1126_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1125 N_OUT9_Mn9@1125_d N_OUT8_Mn9@1125_g N_VSS_Mn9@1125_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1124 N_OUT9_Mn9@1124_d N_OUT8_Mn9@1124_g N_VSS_Mn9@1124_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1125 N_OUT9_Mp9@1125_d N_OUT8_Mp9@1125_g N_VDD_Mp9@1125_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1124 N_OUT9_Mp9@1124_d N_OUT8_Mp9@1124_g N_VDD_Mp9@1124_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1123 N_OUT9_Mn9@1123_d N_OUT8_Mn9@1123_g N_VSS_Mn9@1123_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1122 N_OUT9_Mn9@1122_d N_OUT8_Mn9@1122_g N_VSS_Mn9@1122_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1123 N_OUT9_Mp9@1123_d N_OUT8_Mp9@1123_g N_VDD_Mp9@1123_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1122 N_OUT9_Mp9@1122_d N_OUT8_Mp9@1122_g N_VDD_Mp9@1122_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1121 N_OUT9_Mn9@1121_d N_OUT8_Mn9@1121_g N_VSS_Mn9@1121_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1120 N_OUT9_Mn9@1120_d N_OUT8_Mn9@1120_g N_VSS_Mn9@1120_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1121 N_OUT9_Mp9@1121_d N_OUT8_Mp9@1121_g N_VDD_Mp9@1121_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1120 N_OUT9_Mp9@1120_d N_OUT8_Mp9@1120_g N_VDD_Mp9@1120_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1119 N_OUT9_Mn9@1119_d N_OUT8_Mn9@1119_g N_VSS_Mn9@1119_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1118 N_OUT9_Mn9@1118_d N_OUT8_Mn9@1118_g N_VSS_Mn9@1118_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1119 N_OUT9_Mp9@1119_d N_OUT8_Mp9@1119_g N_VDD_Mp9@1119_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1118 N_OUT9_Mp9@1118_d N_OUT8_Mp9@1118_g N_VDD_Mp9@1118_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1117 N_OUT9_Mn9@1117_d N_OUT8_Mn9@1117_g N_VSS_Mn9@1117_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1116 N_OUT9_Mn9@1116_d N_OUT8_Mn9@1116_g N_VSS_Mn9@1116_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1117 N_OUT9_Mp9@1117_d N_OUT8_Mp9@1117_g N_VDD_Mp9@1117_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1116 N_OUT9_Mp9@1116_d N_OUT8_Mp9@1116_g N_VDD_Mp9@1116_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1115 N_OUT9_Mn9@1115_d N_OUT8_Mn9@1115_g N_VSS_Mn9@1115_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1114 N_OUT9_Mn9@1114_d N_OUT8_Mn9@1114_g N_VSS_Mn9@1114_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1115 N_OUT9_Mp9@1115_d N_OUT8_Mp9@1115_g N_VDD_Mp9@1115_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1114 N_OUT9_Mp9@1114_d N_OUT8_Mp9@1114_g N_VDD_Mp9@1114_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1113 N_OUT9_Mn9@1113_d N_OUT8_Mn9@1113_g N_VSS_Mn9@1113_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1112 N_OUT9_Mn9@1112_d N_OUT8_Mn9@1112_g N_VSS_Mn9@1112_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1113 N_OUT9_Mp9@1113_d N_OUT8_Mp9@1113_g N_VDD_Mp9@1113_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1112 N_OUT9_Mp9@1112_d N_OUT8_Mp9@1112_g N_VDD_Mp9@1112_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1111 N_OUT9_Mn9@1111_d N_OUT8_Mn9@1111_g N_VSS_Mn9@1111_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1110 N_OUT9_Mn9@1110_d N_OUT8_Mn9@1110_g N_VSS_Mn9@1110_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1111 N_OUT9_Mp9@1111_d N_OUT8_Mp9@1111_g N_VDD_Mp9@1111_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1110 N_OUT9_Mp9@1110_d N_OUT8_Mp9@1110_g N_VDD_Mp9@1110_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1109 N_OUT9_Mn9@1109_d N_OUT8_Mn9@1109_g N_VSS_Mn9@1109_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1108 N_OUT9_Mn9@1108_d N_OUT8_Mn9@1108_g N_VSS_Mn9@1108_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1109 N_OUT9_Mp9@1109_d N_OUT8_Mp9@1109_g N_VDD_Mp9@1109_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1108 N_OUT9_Mp9@1108_d N_OUT8_Mp9@1108_g N_VDD_Mp9@1108_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1107 N_OUT9_Mn9@1107_d N_OUT8_Mn9@1107_g N_VSS_Mn9@1107_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1106 N_OUT9_Mn9@1106_d N_OUT8_Mn9@1106_g N_VSS_Mn9@1106_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1107 N_OUT9_Mp9@1107_d N_OUT8_Mp9@1107_g N_VDD_Mp9@1107_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1106 N_OUT9_Mp9@1106_d N_OUT8_Mp9@1106_g N_VDD_Mp9@1106_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1105 N_OUT9_Mn9@1105_d N_OUT8_Mn9@1105_g N_VSS_Mn9@1105_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1104 N_OUT9_Mn9@1104_d N_OUT8_Mn9@1104_g N_VSS_Mn9@1104_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1105 N_OUT9_Mp9@1105_d N_OUT8_Mp9@1105_g N_VDD_Mp9@1105_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1104 N_OUT9_Mp9@1104_d N_OUT8_Mp9@1104_g N_VDD_Mp9@1104_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1103 N_OUT9_Mn9@1103_d N_OUT8_Mn9@1103_g N_VSS_Mn9@1103_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1102 N_OUT9_Mn9@1102_d N_OUT8_Mn9@1102_g N_VSS_Mn9@1102_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1103 N_OUT9_Mp9@1103_d N_OUT8_Mp9@1103_g N_VDD_Mp9@1103_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1102 N_OUT9_Mp9@1102_d N_OUT8_Mp9@1102_g N_VDD_Mp9@1102_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1101 N_OUT9_Mn9@1101_d N_OUT8_Mn9@1101_g N_VSS_Mn9@1101_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1100 N_OUT9_Mn9@1100_d N_OUT8_Mn9@1100_g N_VSS_Mn9@1100_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1101 N_OUT9_Mp9@1101_d N_OUT8_Mp9@1101_g N_VDD_Mp9@1101_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1100 N_OUT9_Mp9@1100_d N_OUT8_Mp9@1100_g N_VDD_Mp9@1100_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1099 N_OUT9_Mn9@1099_d N_OUT8_Mn9@1099_g N_VSS_Mn9@1099_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1098 N_OUT9_Mn9@1098_d N_OUT8_Mn9@1098_g N_VSS_Mn9@1098_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1099 N_OUT9_Mp9@1099_d N_OUT8_Mp9@1099_g N_VDD_Mp9@1099_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1098 N_OUT9_Mp9@1098_d N_OUT8_Mp9@1098_g N_VDD_Mp9@1098_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1097 N_OUT9_Mn9@1097_d N_OUT8_Mn9@1097_g N_VSS_Mn9@1097_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1096 N_OUT9_Mn9@1096_d N_OUT8_Mn9@1096_g N_VSS_Mn9@1096_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1097 N_OUT9_Mp9@1097_d N_OUT8_Mp9@1097_g N_VDD_Mp9@1097_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1096 N_OUT9_Mp9@1096_d N_OUT8_Mp9@1096_g N_VDD_Mp9@1096_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1095 N_OUT9_Mn9@1095_d N_OUT8_Mn9@1095_g N_VSS_Mn9@1095_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1094 N_OUT9_Mn9@1094_d N_OUT8_Mn9@1094_g N_VSS_Mn9@1094_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1095 N_OUT9_Mp9@1095_d N_OUT8_Mp9@1095_g N_VDD_Mp9@1095_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1094 N_OUT9_Mp9@1094_d N_OUT8_Mp9@1094_g N_VDD_Mp9@1094_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1093 N_OUT9_Mn9@1093_d N_OUT8_Mn9@1093_g N_VSS_Mn9@1093_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1092 N_OUT9_Mn9@1092_d N_OUT8_Mn9@1092_g N_VSS_Mn9@1092_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1093 N_OUT9_Mp9@1093_d N_OUT8_Mp9@1093_g N_VDD_Mp9@1093_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1092 N_OUT9_Mp9@1092_d N_OUT8_Mp9@1092_g N_VDD_Mp9@1092_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1091 N_OUT9_Mn9@1091_d N_OUT8_Mn9@1091_g N_VSS_Mn9@1091_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1090 N_OUT9_Mn9@1090_d N_OUT8_Mn9@1090_g N_VSS_Mn9@1090_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1091 N_OUT9_Mp9@1091_d N_OUT8_Mp9@1091_g N_VDD_Mp9@1091_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1090 N_OUT9_Mp9@1090_d N_OUT8_Mp9@1090_g N_VDD_Mp9@1090_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1089 N_OUT9_Mn9@1089_d N_OUT8_Mn9@1089_g N_VSS_Mn9@1089_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1088 N_OUT9_Mn9@1088_d N_OUT8_Mn9@1088_g N_VSS_Mn9@1088_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1089 N_OUT9_Mp9@1089_d N_OUT8_Mp9@1089_g N_VDD_Mp9@1089_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1088 N_OUT9_Mp9@1088_d N_OUT8_Mp9@1088_g N_VDD_Mp9@1088_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1087 N_OUT9_Mn9@1087_d N_OUT8_Mn9@1087_g N_VSS_Mn9@1087_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1086 N_OUT9_Mn9@1086_d N_OUT8_Mn9@1086_g N_VSS_Mn9@1086_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1087 N_OUT9_Mp9@1087_d N_OUT8_Mp9@1087_g N_VDD_Mp9@1087_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1086 N_OUT9_Mp9@1086_d N_OUT8_Mp9@1086_g N_VDD_Mp9@1086_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1085 N_OUT9_Mn9@1085_d N_OUT8_Mn9@1085_g N_VSS_Mn9@1085_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1084 N_OUT9_Mn9@1084_d N_OUT8_Mn9@1084_g N_VSS_Mn9@1084_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1085 N_OUT9_Mp9@1085_d N_OUT8_Mp9@1085_g N_VDD_Mp9@1085_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1084 N_OUT9_Mp9@1084_d N_OUT8_Mp9@1084_g N_VDD_Mp9@1084_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1083 N_OUT9_Mn9@1083_d N_OUT8_Mn9@1083_g N_VSS_Mn9@1083_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1082 N_OUT9_Mn9@1082_d N_OUT8_Mn9@1082_g N_VSS_Mn9@1082_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1083 N_OUT9_Mp9@1083_d N_OUT8_Mp9@1083_g N_VDD_Mp9@1083_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1082 N_OUT9_Mp9@1082_d N_OUT8_Mp9@1082_g N_VDD_Mp9@1082_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1081 N_OUT9_Mn9@1081_d N_OUT8_Mn9@1081_g N_VSS_Mn9@1081_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1080 N_OUT9_Mn9@1080_d N_OUT8_Mn9@1080_g N_VSS_Mn9@1080_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1081 N_OUT9_Mp9@1081_d N_OUT8_Mp9@1081_g N_VDD_Mp9@1081_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1080 N_OUT9_Mp9@1080_d N_OUT8_Mp9@1080_g N_VDD_Mp9@1080_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1079 N_OUT9_Mn9@1079_d N_OUT8_Mn9@1079_g N_VSS_Mn9@1079_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1078 N_OUT9_Mn9@1078_d N_OUT8_Mn9@1078_g N_VSS_Mn9@1078_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1079 N_OUT9_Mp9@1079_d N_OUT8_Mp9@1079_g N_VDD_Mp9@1079_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1078 N_OUT9_Mp9@1078_d N_OUT8_Mp9@1078_g N_VDD_Mp9@1078_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1077 N_OUT9_Mn9@1077_d N_OUT8_Mn9@1077_g N_VSS_Mn9@1077_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1076 N_OUT9_Mn9@1076_d N_OUT8_Mn9@1076_g N_VSS_Mn9@1076_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1077 N_OUT9_Mp9@1077_d N_OUT8_Mp9@1077_g N_VDD_Mp9@1077_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1076 N_OUT9_Mp9@1076_d N_OUT8_Mp9@1076_g N_VDD_Mp9@1076_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1075 N_OUT9_Mn9@1075_d N_OUT8_Mn9@1075_g N_VSS_Mn9@1075_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1074 N_OUT9_Mn9@1074_d N_OUT8_Mn9@1074_g N_VSS_Mn9@1074_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1075 N_OUT9_Mp9@1075_d N_OUT8_Mp9@1075_g N_VDD_Mp9@1075_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1074 N_OUT9_Mp9@1074_d N_OUT8_Mp9@1074_g N_VDD_Mp9@1074_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1073 N_OUT9_Mn9@1073_d N_OUT8_Mn9@1073_g N_VSS_Mn9@1073_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1072 N_OUT9_Mn9@1072_d N_OUT8_Mn9@1072_g N_VSS_Mn9@1072_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1073 N_OUT9_Mp9@1073_d N_OUT8_Mp9@1073_g N_VDD_Mp9@1073_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1072 N_OUT9_Mp9@1072_d N_OUT8_Mp9@1072_g N_VDD_Mp9@1072_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1071 N_OUT9_Mn9@1071_d N_OUT8_Mn9@1071_g N_VSS_Mn9@1071_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1070 N_OUT9_Mn9@1070_d N_OUT8_Mn9@1070_g N_VSS_Mn9@1070_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1071 N_OUT9_Mp9@1071_d N_OUT8_Mp9@1071_g N_VDD_Mp9@1071_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1070 N_OUT9_Mp9@1070_d N_OUT8_Mp9@1070_g N_VDD_Mp9@1070_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1069 N_OUT9_Mn9@1069_d N_OUT8_Mn9@1069_g N_VSS_Mn9@1069_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1068 N_OUT9_Mn9@1068_d N_OUT8_Mn9@1068_g N_VSS_Mn9@1068_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1069 N_OUT9_Mp9@1069_d N_OUT8_Mp9@1069_g N_VDD_Mp9@1069_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1068 N_OUT9_Mp9@1068_d N_OUT8_Mp9@1068_g N_VDD_Mp9@1068_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1067 N_OUT9_Mn9@1067_d N_OUT8_Mn9@1067_g N_VSS_Mn9@1067_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1066 N_OUT9_Mn9@1066_d N_OUT8_Mn9@1066_g N_VSS_Mn9@1066_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1067 N_OUT9_Mp9@1067_d N_OUT8_Mp9@1067_g N_VDD_Mp9@1067_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1066 N_OUT9_Mp9@1066_d N_OUT8_Mp9@1066_g N_VDD_Mp9@1066_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1065 N_OUT9_Mn9@1065_d N_OUT8_Mn9@1065_g N_VSS_Mn9@1065_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1064 N_OUT9_Mn9@1064_d N_OUT8_Mn9@1064_g N_VSS_Mn9@1064_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1065 N_OUT9_Mp9@1065_d N_OUT8_Mp9@1065_g N_VDD_Mp9@1065_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1064 N_OUT9_Mp9@1064_d N_OUT8_Mp9@1064_g N_VDD_Mp9@1064_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1063 N_OUT9_Mn9@1063_d N_OUT8_Mn9@1063_g N_VSS_Mn9@1063_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1062 N_OUT9_Mn9@1062_d N_OUT8_Mn9@1062_g N_VSS_Mn9@1062_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1063 N_OUT9_Mp9@1063_d N_OUT8_Mp9@1063_g N_VDD_Mp9@1063_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1062 N_OUT9_Mp9@1062_d N_OUT8_Mp9@1062_g N_VDD_Mp9@1062_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1061 N_OUT9_Mn9@1061_d N_OUT8_Mn9@1061_g N_VSS_Mn9@1061_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1060 N_OUT9_Mn9@1060_d N_OUT8_Mn9@1060_g N_VSS_Mn9@1060_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1061 N_OUT9_Mp9@1061_d N_OUT8_Mp9@1061_g N_VDD_Mp9@1061_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1060 N_OUT9_Mp9@1060_d N_OUT8_Mp9@1060_g N_VDD_Mp9@1060_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1059 N_OUT9_Mn9@1059_d N_OUT8_Mn9@1059_g N_VSS_Mn9@1059_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1058 N_OUT9_Mn9@1058_d N_OUT8_Mn9@1058_g N_VSS_Mn9@1058_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1059 N_OUT9_Mp9@1059_d N_OUT8_Mp9@1059_g N_VDD_Mp9@1059_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1058 N_OUT9_Mp9@1058_d N_OUT8_Mp9@1058_g N_VDD_Mp9@1058_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1057 N_OUT9_Mn9@1057_d N_OUT8_Mn9@1057_g N_VSS_Mn9@1057_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1056 N_OUT9_Mn9@1056_d N_OUT8_Mn9@1056_g N_VSS_Mn9@1056_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1057 N_OUT9_Mp9@1057_d N_OUT8_Mp9@1057_g N_VDD_Mp9@1057_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1056 N_OUT9_Mp9@1056_d N_OUT8_Mp9@1056_g N_VDD_Mp9@1056_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1055 N_OUT9_Mn9@1055_d N_OUT8_Mn9@1055_g N_VSS_Mn9@1055_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1054 N_OUT9_Mn9@1054_d N_OUT8_Mn9@1054_g N_VSS_Mn9@1054_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1055 N_OUT9_Mp9@1055_d N_OUT8_Mp9@1055_g N_VDD_Mp9@1055_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1054 N_OUT9_Mp9@1054_d N_OUT8_Mp9@1054_g N_VDD_Mp9@1054_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1053 N_OUT9_Mn9@1053_d N_OUT8_Mn9@1053_g N_VSS_Mn9@1053_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1052 N_OUT9_Mn9@1052_d N_OUT8_Mn9@1052_g N_VSS_Mn9@1052_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1053 N_OUT9_Mp9@1053_d N_OUT8_Mp9@1053_g N_VDD_Mp9@1053_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1052 N_OUT9_Mp9@1052_d N_OUT8_Mp9@1052_g N_VDD_Mp9@1052_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1051 N_OUT9_Mn9@1051_d N_OUT8_Mn9@1051_g N_VSS_Mn9@1051_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1050 N_OUT9_Mn9@1050_d N_OUT8_Mn9@1050_g N_VSS_Mn9@1050_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1051 N_OUT9_Mp9@1051_d N_OUT8_Mp9@1051_g N_VDD_Mp9@1051_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1050 N_OUT9_Mp9@1050_d N_OUT8_Mp9@1050_g N_VDD_Mp9@1050_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1049 N_OUT9_Mn9@1049_d N_OUT8_Mn9@1049_g N_VSS_Mn9@1049_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1048 N_OUT9_Mn9@1048_d N_OUT8_Mn9@1048_g N_VSS_Mn9@1048_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1049 N_OUT9_Mp9@1049_d N_OUT8_Mp9@1049_g N_VDD_Mp9@1049_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1048 N_OUT9_Mp9@1048_d N_OUT8_Mp9@1048_g N_VDD_Mp9@1048_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1047 N_OUT9_Mn9@1047_d N_OUT8_Mn9@1047_g N_VSS_Mn9@1047_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1046 N_OUT9_Mn9@1046_d N_OUT8_Mn9@1046_g N_VSS_Mn9@1046_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1047 N_OUT9_Mp9@1047_d N_OUT8_Mp9@1047_g N_VDD_Mp9@1047_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1046 N_OUT9_Mp9@1046_d N_OUT8_Mp9@1046_g N_VDD_Mp9@1046_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1045 N_OUT9_Mn9@1045_d N_OUT8_Mn9@1045_g N_VSS_Mn9@1045_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1044 N_OUT9_Mn9@1044_d N_OUT8_Mn9@1044_g N_VSS_Mn9@1044_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1045 N_OUT9_Mp9@1045_d N_OUT8_Mp9@1045_g N_VDD_Mp9@1045_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1044 N_OUT9_Mp9@1044_d N_OUT8_Mp9@1044_g N_VDD_Mp9@1044_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1043 N_OUT9_Mn9@1043_d N_OUT8_Mn9@1043_g N_VSS_Mn9@1043_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1042 N_OUT9_Mn9@1042_d N_OUT8_Mn9@1042_g N_VSS_Mn9@1042_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1043 N_OUT9_Mp9@1043_d N_OUT8_Mp9@1043_g N_VDD_Mp9@1043_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1042 N_OUT9_Mp9@1042_d N_OUT8_Mp9@1042_g N_VDD_Mp9@1042_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1041 N_OUT9_Mn9@1041_d N_OUT8_Mn9@1041_g N_VSS_Mn9@1041_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1040 N_OUT9_Mn9@1040_d N_OUT8_Mn9@1040_g N_VSS_Mn9@1040_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1041 N_OUT9_Mp9@1041_d N_OUT8_Mp9@1041_g N_VDD_Mp9@1041_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1040 N_OUT9_Mp9@1040_d N_OUT8_Mp9@1040_g N_VDD_Mp9@1040_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1039 N_OUT9_Mn9@1039_d N_OUT8_Mn9@1039_g N_VSS_Mn9@1039_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1038 N_OUT9_Mn9@1038_d N_OUT8_Mn9@1038_g N_VSS_Mn9@1038_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1039 N_OUT9_Mp9@1039_d N_OUT8_Mp9@1039_g N_VDD_Mp9@1039_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1038 N_OUT9_Mp9@1038_d N_OUT8_Mp9@1038_g N_VDD_Mp9@1038_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1037 N_OUT9_Mn9@1037_d N_OUT8_Mn9@1037_g N_VSS_Mn9@1037_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1036 N_OUT9_Mn9@1036_d N_OUT8_Mn9@1036_g N_VSS_Mn9@1036_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1037 N_OUT9_Mp9@1037_d N_OUT8_Mp9@1037_g N_VDD_Mp9@1037_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1036 N_OUT9_Mp9@1036_d N_OUT8_Mp9@1036_g N_VDD_Mp9@1036_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1035 N_OUT9_Mn9@1035_d N_OUT8_Mn9@1035_g N_VSS_Mn9@1035_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1034 N_OUT9_Mn9@1034_d N_OUT8_Mn9@1034_g N_VSS_Mn9@1034_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1035 N_OUT9_Mp9@1035_d N_OUT8_Mp9@1035_g N_VDD_Mp9@1035_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1034 N_OUT9_Mp9@1034_d N_OUT8_Mp9@1034_g N_VDD_Mp9@1034_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1033 N_OUT9_Mn9@1033_d N_OUT8_Mn9@1033_g N_VSS_Mn9@1033_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1032 N_OUT9_Mn9@1032_d N_OUT8_Mn9@1032_g N_VSS_Mn9@1032_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1033 N_OUT9_Mp9@1033_d N_OUT8_Mp9@1033_g N_VDD_Mp9@1033_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1032 N_OUT9_Mp9@1032_d N_OUT8_Mp9@1032_g N_VDD_Mp9@1032_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1031 N_OUT9_Mn9@1031_d N_OUT8_Mn9@1031_g N_VSS_Mn9@1031_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1030 N_OUT9_Mn9@1030_d N_OUT8_Mn9@1030_g N_VSS_Mn9@1030_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1031 N_OUT9_Mp9@1031_d N_OUT8_Mp9@1031_g N_VDD_Mp9@1031_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1030 N_OUT9_Mp9@1030_d N_OUT8_Mp9@1030_g N_VDD_Mp9@1030_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1029 N_OUT9_Mn9@1029_d N_OUT8_Mn9@1029_g N_VSS_Mn9@1029_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1028 N_OUT9_Mn9@1028_d N_OUT8_Mn9@1028_g N_VSS_Mn9@1028_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1029 N_OUT9_Mp9@1029_d N_OUT8_Mp9@1029_g N_VDD_Mp9@1029_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1028 N_OUT9_Mp9@1028_d N_OUT8_Mp9@1028_g N_VDD_Mp9@1028_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1027 N_OUT9_Mn9@1027_d N_OUT8_Mn9@1027_g N_VSS_Mn9@1027_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1026 N_OUT9_Mn9@1026_d N_OUT8_Mn9@1026_g N_VSS_Mn9@1026_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1027 N_OUT9_Mp9@1027_d N_OUT8_Mp9@1027_g N_VDD_Mp9@1027_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1026 N_OUT9_Mp9@1026_d N_OUT8_Mp9@1026_g N_VDD_Mp9@1026_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1025 N_OUT9_Mn9@1025_d N_OUT8_Mn9@1025_g N_VSS_Mn9@1025_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1024 N_OUT9_Mn9@1024_d N_OUT8_Mn9@1024_g N_VSS_Mn9@1024_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1025 N_OUT9_Mp9@1025_d N_OUT8_Mp9@1025_g N_VDD_Mp9@1025_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1024 N_OUT9_Mp9@1024_d N_OUT8_Mp9@1024_g N_VDD_Mp9@1024_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1023 N_OUT9_Mn9@1023_d N_OUT8_Mn9@1023_g N_VSS_Mn9@1023_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1022 N_OUT9_Mn9@1022_d N_OUT8_Mn9@1022_g N_VSS_Mn9@1022_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1023 N_OUT9_Mp9@1023_d N_OUT8_Mp9@1023_g N_VDD_Mp9@1023_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1022 N_OUT9_Mp9@1022_d N_OUT8_Mp9@1022_g N_VDD_Mp9@1022_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1021 N_OUT9_Mn9@1021_d N_OUT8_Mn9@1021_g N_VSS_Mn9@1021_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1020 N_OUT9_Mn9@1020_d N_OUT8_Mn9@1020_g N_VSS_Mn9@1020_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1021 N_OUT9_Mp9@1021_d N_OUT8_Mp9@1021_g N_VDD_Mp9@1021_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1020 N_OUT9_Mp9@1020_d N_OUT8_Mp9@1020_g N_VDD_Mp9@1020_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1019 N_OUT9_Mn9@1019_d N_OUT8_Mn9@1019_g N_VSS_Mn9@1019_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1018 N_OUT9_Mn9@1018_d N_OUT8_Mn9@1018_g N_VSS_Mn9@1018_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1019 N_OUT9_Mp9@1019_d N_OUT8_Mp9@1019_g N_VDD_Mp9@1019_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1018 N_OUT9_Mp9@1018_d N_OUT8_Mp9@1018_g N_VDD_Mp9@1018_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1017 N_OUT9_Mn9@1017_d N_OUT8_Mn9@1017_g N_VSS_Mn9@1017_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1016 N_OUT9_Mn9@1016_d N_OUT8_Mn9@1016_g N_VSS_Mn9@1016_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1017 N_OUT9_Mp9@1017_d N_OUT8_Mp9@1017_g N_VDD_Mp9@1017_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1016 N_OUT9_Mp9@1016_d N_OUT8_Mp9@1016_g N_VDD_Mp9@1016_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1015 N_OUT9_Mn9@1015_d N_OUT8_Mn9@1015_g N_VSS_Mn9@1015_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1014 N_OUT9_Mn9@1014_d N_OUT8_Mn9@1014_g N_VSS_Mn9@1014_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1015 N_OUT9_Mp9@1015_d N_OUT8_Mp9@1015_g N_VDD_Mp9@1015_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1014 N_OUT9_Mp9@1014_d N_OUT8_Mp9@1014_g N_VDD_Mp9@1014_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1013 N_OUT9_Mn9@1013_d N_OUT8_Mn9@1013_g N_VSS_Mn9@1013_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1012 N_OUT9_Mn9@1012_d N_OUT8_Mn9@1012_g N_VSS_Mn9@1012_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1013 N_OUT9_Mp9@1013_d N_OUT8_Mp9@1013_g N_VDD_Mp9@1013_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1012 N_OUT9_Mp9@1012_d N_OUT8_Mp9@1012_g N_VDD_Mp9@1012_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1011 N_OUT9_Mn9@1011_d N_OUT8_Mn9@1011_g N_VSS_Mn9@1011_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1010 N_OUT9_Mn9@1010_d N_OUT8_Mn9@1010_g N_VSS_Mn9@1010_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1011 N_OUT9_Mp9@1011_d N_OUT8_Mp9@1011_g N_VDD_Mp9@1011_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1010 N_OUT9_Mp9@1010_d N_OUT8_Mp9@1010_g N_VDD_Mp9@1010_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1009 N_OUT9_Mn9@1009_d N_OUT8_Mn9@1009_g N_VSS_Mn9@1009_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1008 N_OUT9_Mn9@1008_d N_OUT8_Mn9@1008_g N_VSS_Mn9@1008_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1009 N_OUT9_Mp9@1009_d N_OUT8_Mp9@1009_g N_VDD_Mp9@1009_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1008 N_OUT9_Mp9@1008_d N_OUT8_Mp9@1008_g N_VDD_Mp9@1008_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1007 N_OUT9_Mn9@1007_d N_OUT8_Mn9@1007_g N_VSS_Mn9@1007_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1006 N_OUT9_Mn9@1006_d N_OUT8_Mn9@1006_g N_VSS_Mn9@1006_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1007 N_OUT9_Mp9@1007_d N_OUT8_Mp9@1007_g N_VDD_Mp9@1007_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1006 N_OUT9_Mp9@1006_d N_OUT8_Mp9@1006_g N_VDD_Mp9@1006_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1005 N_OUT9_Mn9@1005_d N_OUT8_Mn9@1005_g N_VSS_Mn9@1005_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1004 N_OUT9_Mn9@1004_d N_OUT8_Mn9@1004_g N_VSS_Mn9@1004_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1005 N_OUT9_Mp9@1005_d N_OUT8_Mp9@1005_g N_VDD_Mp9@1005_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1004 N_OUT9_Mp9@1004_d N_OUT8_Mp9@1004_g N_VDD_Mp9@1004_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1003 N_OUT9_Mn9@1003_d N_OUT8_Mn9@1003_g N_VSS_Mn9@1003_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1002 N_OUT9_Mn9@1002_d N_OUT8_Mn9@1002_g N_VSS_Mn9@1002_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1003 N_OUT9_Mp9@1003_d N_OUT8_Mp9@1003_g N_VDD_Mp9@1003_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1002 N_OUT9_Mp9@1002_d N_OUT8_Mp9@1002_g N_VDD_Mp9@1002_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@1001 N_OUT9_Mn9@1001_d N_OUT8_Mn9@1001_g N_VSS_Mn9@1001_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@1000 N_OUT9_Mn9@1000_d N_OUT8_Mn9@1000_g N_VSS_Mn9@1000_s N_VSS_Mn7@1159_b
+ N_18 L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@1001 N_OUT9_Mp9@1001_d N_OUT8_Mp9@1001_g N_VDD_Mp9@1001_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@1000 N_OUT9_Mp9@1000_d N_OUT8_Mp9@1000_g N_VDD_Mp9@1000_s N_VDD_Mp9@4995_b
+ P_18 L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@999 N_OUT9_Mn9@999_d N_OUT8_Mn9@999_g N_VSS_Mn9@999_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@998 N_OUT9_Mn9@998_d N_OUT8_Mn9@998_g N_VSS_Mn9@998_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@999 N_OUT9_Mp9@999_d N_OUT8_Mp9@999_g N_VDD_Mp9@999_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@998 N_OUT9_Mp9@998_d N_OUT8_Mp9@998_g N_VDD_Mp9@998_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@997 N_OUT9_Mn9@997_d N_OUT8_Mn9@997_g N_VSS_Mn9@997_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@996 N_OUT9_Mn9@996_d N_OUT8_Mn9@996_g N_VSS_Mn9@996_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@997 N_OUT9_Mp9@997_d N_OUT8_Mp9@997_g N_VDD_Mp9@997_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@996 N_OUT9_Mp9@996_d N_OUT8_Mp9@996_g N_VDD_Mp9@996_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@995 N_OUT9_Mn9@995_d N_OUT8_Mn9@995_g N_VSS_Mn9@995_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@994 N_OUT9_Mn9@994_d N_OUT8_Mn9@994_g N_VSS_Mn9@994_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@995 N_OUT9_Mp9@995_d N_OUT8_Mp9@995_g N_VDD_Mp9@995_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@994 N_OUT9_Mp9@994_d N_OUT8_Mp9@994_g N_VDD_Mp9@994_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@993 N_OUT9_Mn9@993_d N_OUT8_Mn9@993_g N_VSS_Mn9@993_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@992 N_OUT9_Mn9@992_d N_OUT8_Mn9@992_g N_VSS_Mn9@992_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@993 N_OUT9_Mp9@993_d N_OUT8_Mp9@993_g N_VDD_Mp9@993_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@992 N_OUT9_Mp9@992_d N_OUT8_Mp9@992_g N_VDD_Mp9@992_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@991 N_OUT9_Mn9@991_d N_OUT8_Mn9@991_g N_VSS_Mn9@991_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@990 N_OUT9_Mn9@990_d N_OUT8_Mn9@990_g N_VSS_Mn9@990_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@991 N_OUT9_Mp9@991_d N_OUT8_Mp9@991_g N_VDD_Mp9@991_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@990 N_OUT9_Mp9@990_d N_OUT8_Mp9@990_g N_VDD_Mp9@990_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@989 N_OUT9_Mn9@989_d N_OUT8_Mn9@989_g N_VSS_Mn9@989_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@988 N_OUT9_Mn9@988_d N_OUT8_Mn9@988_g N_VSS_Mn9@988_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@989 N_OUT9_Mp9@989_d N_OUT8_Mp9@989_g N_VDD_Mp9@989_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@988 N_OUT9_Mp9@988_d N_OUT8_Mp9@988_g N_VDD_Mp9@988_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@987 N_OUT9_Mn9@987_d N_OUT8_Mn9@987_g N_VSS_Mn9@987_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@986 N_OUT9_Mn9@986_d N_OUT8_Mn9@986_g N_VSS_Mn9@986_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@987 N_OUT9_Mp9@987_d N_OUT8_Mp9@987_g N_VDD_Mp9@987_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@986 N_OUT9_Mp9@986_d N_OUT8_Mp9@986_g N_VDD_Mp9@986_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@985 N_OUT9_Mn9@985_d N_OUT8_Mn9@985_g N_VSS_Mn9@985_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@984 N_OUT9_Mn9@984_d N_OUT8_Mn9@984_g N_VSS_Mn9@984_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@985 N_OUT9_Mp9@985_d N_OUT8_Mp9@985_g N_VDD_Mp9@985_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@984 N_OUT9_Mp9@984_d N_OUT8_Mp9@984_g N_VDD_Mp9@984_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@983 N_OUT9_Mn9@983_d N_OUT8_Mn9@983_g N_VSS_Mn9@983_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@982 N_OUT9_Mn9@982_d N_OUT8_Mn9@982_g N_VSS_Mn9@982_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@983 N_OUT9_Mp9@983_d N_OUT8_Mp9@983_g N_VDD_Mp9@983_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@982 N_OUT9_Mp9@982_d N_OUT8_Mp9@982_g N_VDD_Mp9@982_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@981 N_OUT9_Mn9@981_d N_OUT8_Mn9@981_g N_VSS_Mn9@981_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@980 N_OUT9_Mn9@980_d N_OUT8_Mn9@980_g N_VSS_Mn9@980_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@981 N_OUT9_Mp9@981_d N_OUT8_Mp9@981_g N_VDD_Mp9@981_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@980 N_OUT9_Mp9@980_d N_OUT8_Mp9@980_g N_VDD_Mp9@980_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@979 N_OUT9_Mn9@979_d N_OUT8_Mn9@979_g N_VSS_Mn9@979_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@978 N_OUT9_Mn9@978_d N_OUT8_Mn9@978_g N_VSS_Mn9@978_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@979 N_OUT9_Mp9@979_d N_OUT8_Mp9@979_g N_VDD_Mp9@979_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@978 N_OUT9_Mp9@978_d N_OUT8_Mp9@978_g N_VDD_Mp9@978_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@977 N_OUT9_Mn9@977_d N_OUT8_Mn9@977_g N_VSS_Mn9@977_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@976 N_OUT9_Mn9@976_d N_OUT8_Mn9@976_g N_VSS_Mn9@976_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@977 N_OUT9_Mp9@977_d N_OUT8_Mp9@977_g N_VDD_Mp9@977_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@976 N_OUT9_Mp9@976_d N_OUT8_Mp9@976_g N_VDD_Mp9@976_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@975 N_OUT9_Mn9@975_d N_OUT8_Mn9@975_g N_VSS_Mn9@975_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@974 N_OUT9_Mn9@974_d N_OUT8_Mn9@974_g N_VSS_Mn9@974_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@975 N_OUT9_Mp9@975_d N_OUT8_Mp9@975_g N_VDD_Mp9@975_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@974 N_OUT9_Mp9@974_d N_OUT8_Mp9@974_g N_VDD_Mp9@974_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@973 N_OUT9_Mn9@973_d N_OUT8_Mn9@973_g N_VSS_Mn9@973_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@972 N_OUT9_Mn9@972_d N_OUT8_Mn9@972_g N_VSS_Mn9@972_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@973 N_OUT9_Mp9@973_d N_OUT8_Mp9@973_g N_VDD_Mp9@973_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@972 N_OUT9_Mp9@972_d N_OUT8_Mp9@972_g N_VDD_Mp9@972_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@971 N_OUT9_Mn9@971_d N_OUT8_Mn9@971_g N_VSS_Mn9@971_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@970 N_OUT9_Mn9@970_d N_OUT8_Mn9@970_g N_VSS_Mn9@970_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@971 N_OUT9_Mp9@971_d N_OUT8_Mp9@971_g N_VDD_Mp9@971_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@970 N_OUT9_Mp9@970_d N_OUT8_Mp9@970_g N_VDD_Mp9@970_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@969 N_OUT9_Mn9@969_d N_OUT8_Mn9@969_g N_VSS_Mn9@969_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@968 N_OUT9_Mn9@968_d N_OUT8_Mn9@968_g N_VSS_Mn9@968_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@969 N_OUT9_Mp9@969_d N_OUT8_Mp9@969_g N_VDD_Mp9@969_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@968 N_OUT9_Mp9@968_d N_OUT8_Mp9@968_g N_VDD_Mp9@968_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@967 N_OUT9_Mn9@967_d N_OUT8_Mn9@967_g N_VSS_Mn9@967_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@966 N_OUT9_Mn9@966_d N_OUT8_Mn9@966_g N_VSS_Mn9@966_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@967 N_OUT9_Mp9@967_d N_OUT8_Mp9@967_g N_VDD_Mp9@967_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@966 N_OUT9_Mp9@966_d N_OUT8_Mp9@966_g N_VDD_Mp9@966_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@965 N_OUT9_Mn9@965_d N_OUT8_Mn9@965_g N_VSS_Mn9@965_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@964 N_OUT9_Mn9@964_d N_OUT8_Mn9@964_g N_VSS_Mn9@964_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@965 N_OUT9_Mp9@965_d N_OUT8_Mp9@965_g N_VDD_Mp9@965_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@964 N_OUT9_Mp9@964_d N_OUT8_Mp9@964_g N_VDD_Mp9@964_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@963 N_OUT9_Mn9@963_d N_OUT8_Mn9@963_g N_VSS_Mn9@963_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@962 N_OUT9_Mn9@962_d N_OUT8_Mn9@962_g N_VSS_Mn9@962_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@963 N_OUT9_Mp9@963_d N_OUT8_Mp9@963_g N_VDD_Mp9@963_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@962 N_OUT9_Mp9@962_d N_OUT8_Mp9@962_g N_VDD_Mp9@962_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@961 N_OUT9_Mn9@961_d N_OUT8_Mn9@961_g N_VSS_Mn9@961_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@960 N_OUT9_Mn9@960_d N_OUT8_Mn9@960_g N_VSS_Mn9@960_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@961 N_OUT9_Mp9@961_d N_OUT8_Mp9@961_g N_VDD_Mp9@961_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@960 N_OUT9_Mp9@960_d N_OUT8_Mp9@960_g N_VDD_Mp9@960_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@959 N_OUT9_Mn9@959_d N_OUT8_Mn9@959_g N_VSS_Mn9@959_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@958 N_OUT9_Mn9@958_d N_OUT8_Mn9@958_g N_VSS_Mn9@958_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@959 N_OUT9_Mp9@959_d N_OUT8_Mp9@959_g N_VDD_Mp9@959_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@958 N_OUT9_Mp9@958_d N_OUT8_Mp9@958_g N_VDD_Mp9@958_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@957 N_OUT9_Mn9@957_d N_OUT8_Mn9@957_g N_VSS_Mn9@957_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@956 N_OUT9_Mn9@956_d N_OUT8_Mn9@956_g N_VSS_Mn9@956_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@957 N_OUT9_Mp9@957_d N_OUT8_Mp9@957_g N_VDD_Mp9@957_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@956 N_OUT9_Mp9@956_d N_OUT8_Mp9@956_g N_VDD_Mp9@956_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@955 N_OUT9_Mn9@955_d N_OUT8_Mn9@955_g N_VSS_Mn9@955_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@954 N_OUT9_Mn9@954_d N_OUT8_Mn9@954_g N_VSS_Mn9@954_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@955 N_OUT9_Mp9@955_d N_OUT8_Mp9@955_g N_VDD_Mp9@955_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@954 N_OUT9_Mp9@954_d N_OUT8_Mp9@954_g N_VDD_Mp9@954_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@953 N_OUT9_Mn9@953_d N_OUT8_Mn9@953_g N_VSS_Mn9@953_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@952 N_OUT9_Mn9@952_d N_OUT8_Mn9@952_g N_VSS_Mn9@952_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@953 N_OUT9_Mp9@953_d N_OUT8_Mp9@953_g N_VDD_Mp9@953_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@952 N_OUT9_Mp9@952_d N_OUT8_Mp9@952_g N_VDD_Mp9@952_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@951 N_OUT9_Mn9@951_d N_OUT8_Mn9@951_g N_VSS_Mn9@951_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@950 N_OUT9_Mn9@950_d N_OUT8_Mn9@950_g N_VSS_Mn9@950_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@951 N_OUT9_Mp9@951_d N_OUT8_Mp9@951_g N_VDD_Mp9@951_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@950 N_OUT9_Mp9@950_d N_OUT8_Mp9@950_g N_VDD_Mp9@950_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@949 N_OUT9_Mn9@949_d N_OUT8_Mn9@949_g N_VSS_Mn9@949_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@948 N_OUT9_Mn9@948_d N_OUT8_Mn9@948_g N_VSS_Mn9@948_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@949 N_OUT9_Mp9@949_d N_OUT8_Mp9@949_g N_VDD_Mp9@949_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@948 N_OUT9_Mp9@948_d N_OUT8_Mp9@948_g N_VDD_Mp9@948_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@947 N_OUT9_Mn9@947_d N_OUT8_Mn9@947_g N_VSS_Mn9@947_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@946 N_OUT9_Mn9@946_d N_OUT8_Mn9@946_g N_VSS_Mn9@946_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@947 N_OUT9_Mp9@947_d N_OUT8_Mp9@947_g N_VDD_Mp9@947_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@946 N_OUT9_Mp9@946_d N_OUT8_Mp9@946_g N_VDD_Mp9@946_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@945 N_OUT9_Mn9@945_d N_OUT8_Mn9@945_g N_VSS_Mn9@945_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@944 N_OUT9_Mn9@944_d N_OUT8_Mn9@944_g N_VSS_Mn9@944_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@945 N_OUT9_Mp9@945_d N_OUT8_Mp9@945_g N_VDD_Mp9@945_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@944 N_OUT9_Mp9@944_d N_OUT8_Mp9@944_g N_VDD_Mp9@944_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@943 N_OUT9_Mn9@943_d N_OUT8_Mn9@943_g N_VSS_Mn9@943_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@942 N_OUT9_Mn9@942_d N_OUT8_Mn9@942_g N_VSS_Mn9@942_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@943 N_OUT9_Mp9@943_d N_OUT8_Mp9@943_g N_VDD_Mp9@943_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@942 N_OUT9_Mp9@942_d N_OUT8_Mp9@942_g N_VDD_Mp9@942_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@941 N_OUT9_Mn9@941_d N_OUT8_Mn9@941_g N_VSS_Mn9@941_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@940 N_OUT9_Mn9@940_d N_OUT8_Mn9@940_g N_VSS_Mn9@940_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@941 N_OUT9_Mp9@941_d N_OUT8_Mp9@941_g N_VDD_Mp9@941_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@940 N_OUT9_Mp9@940_d N_OUT8_Mp9@940_g N_VDD_Mp9@940_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@939 N_OUT9_Mn9@939_d N_OUT8_Mn9@939_g N_VSS_Mn9@939_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@938 N_OUT9_Mn9@938_d N_OUT8_Mn9@938_g N_VSS_Mn9@938_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@939 N_OUT9_Mp9@939_d N_OUT8_Mp9@939_g N_VDD_Mp9@939_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@938 N_OUT9_Mp9@938_d N_OUT8_Mp9@938_g N_VDD_Mp9@938_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@937 N_OUT9_Mn9@937_d N_OUT8_Mn9@937_g N_VSS_Mn9@937_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@936 N_OUT9_Mn9@936_d N_OUT8_Mn9@936_g N_VSS_Mn9@936_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@937 N_OUT9_Mp9@937_d N_OUT8_Mp9@937_g N_VDD_Mp9@937_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@936 N_OUT9_Mp9@936_d N_OUT8_Mp9@936_g N_VDD_Mp9@936_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@935 N_OUT9_Mn9@935_d N_OUT8_Mn9@935_g N_VSS_Mn9@935_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@934 N_OUT9_Mn9@934_d N_OUT8_Mn9@934_g N_VSS_Mn9@934_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@935 N_OUT9_Mp9@935_d N_OUT8_Mp9@935_g N_VDD_Mp9@935_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@934 N_OUT9_Mp9@934_d N_OUT8_Mp9@934_g N_VDD_Mp9@934_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@933 N_OUT9_Mn9@933_d N_OUT8_Mn9@933_g N_VSS_Mn9@933_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@932 N_OUT9_Mn9@932_d N_OUT8_Mn9@932_g N_VSS_Mn9@932_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@933 N_OUT9_Mp9@933_d N_OUT8_Mp9@933_g N_VDD_Mp9@933_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@932 N_OUT9_Mp9@932_d N_OUT8_Mp9@932_g N_VDD_Mp9@932_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@931 N_OUT9_Mn9@931_d N_OUT8_Mn9@931_g N_VSS_Mn9@931_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@930 N_OUT9_Mn9@930_d N_OUT8_Mn9@930_g N_VSS_Mn9@930_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@931 N_OUT9_Mp9@931_d N_OUT8_Mp9@931_g N_VDD_Mp9@931_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@930 N_OUT9_Mp9@930_d N_OUT8_Mp9@930_g N_VDD_Mp9@930_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@929 N_OUT9_Mn9@929_d N_OUT8_Mn9@929_g N_VSS_Mn9@929_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@928 N_OUT9_Mn9@928_d N_OUT8_Mn9@928_g N_VSS_Mn9@928_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@929 N_OUT9_Mp9@929_d N_OUT8_Mp9@929_g N_VDD_Mp9@929_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@928 N_OUT9_Mp9@928_d N_OUT8_Mp9@928_g N_VDD_Mp9@928_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@927 N_OUT9_Mn9@927_d N_OUT8_Mn9@927_g N_VSS_Mn9@927_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@926 N_OUT9_Mn9@926_d N_OUT8_Mn9@926_g N_VSS_Mn9@926_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@927 N_OUT9_Mp9@927_d N_OUT8_Mp9@927_g N_VDD_Mp9@927_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@926 N_OUT9_Mp9@926_d N_OUT8_Mp9@926_g N_VDD_Mp9@926_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@925 N_OUT9_Mn9@925_d N_OUT8_Mn9@925_g N_VSS_Mn9@925_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@924 N_OUT9_Mn9@924_d N_OUT8_Mn9@924_g N_VSS_Mn9@924_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@925 N_OUT9_Mp9@925_d N_OUT8_Mp9@925_g N_VDD_Mp9@925_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@924 N_OUT9_Mp9@924_d N_OUT8_Mp9@924_g N_VDD_Mp9@924_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@923 N_OUT9_Mn9@923_d N_OUT8_Mn9@923_g N_VSS_Mn9@923_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@922 N_OUT9_Mn9@922_d N_OUT8_Mn9@922_g N_VSS_Mn9@922_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@923 N_OUT9_Mp9@923_d N_OUT8_Mp9@923_g N_VDD_Mp9@923_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@922 N_OUT9_Mp9@922_d N_OUT8_Mp9@922_g N_VDD_Mp9@922_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@921 N_OUT9_Mn9@921_d N_OUT8_Mn9@921_g N_VSS_Mn9@921_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@920 N_OUT9_Mn9@920_d N_OUT8_Mn9@920_g N_VSS_Mn9@920_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@921 N_OUT9_Mp9@921_d N_OUT8_Mp9@921_g N_VDD_Mp9@921_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@920 N_OUT9_Mp9@920_d N_OUT8_Mp9@920_g N_VDD_Mp9@920_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@919 N_OUT9_Mn9@919_d N_OUT8_Mn9@919_g N_VSS_Mn9@919_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@918 N_OUT9_Mn9@918_d N_OUT8_Mn9@918_g N_VSS_Mn9@918_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@919 N_OUT9_Mp9@919_d N_OUT8_Mp9@919_g N_VDD_Mp9@919_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@918 N_OUT9_Mp9@918_d N_OUT8_Mp9@918_g N_VDD_Mp9@918_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@917 N_OUT9_Mn9@917_d N_OUT8_Mn9@917_g N_VSS_Mn9@917_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@916 N_OUT9_Mn9@916_d N_OUT8_Mn9@916_g N_VSS_Mn9@916_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@917 N_OUT9_Mp9@917_d N_OUT8_Mp9@917_g N_VDD_Mp9@917_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@916 N_OUT9_Mp9@916_d N_OUT8_Mp9@916_g N_VDD_Mp9@916_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@915 N_OUT9_Mn9@915_d N_OUT8_Mn9@915_g N_VSS_Mn9@915_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@914 N_OUT9_Mn9@914_d N_OUT8_Mn9@914_g N_VSS_Mn9@914_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@915 N_OUT9_Mp9@915_d N_OUT8_Mp9@915_g N_VDD_Mp9@915_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@914 N_OUT9_Mp9@914_d N_OUT8_Mp9@914_g N_VDD_Mp9@914_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@913 N_OUT9_Mn9@913_d N_OUT8_Mn9@913_g N_VSS_Mn9@913_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@912 N_OUT9_Mn9@912_d N_OUT8_Mn9@912_g N_VSS_Mn9@912_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@913 N_OUT9_Mp9@913_d N_OUT8_Mp9@913_g N_VDD_Mp9@913_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@912 N_OUT9_Mp9@912_d N_OUT8_Mp9@912_g N_VDD_Mp9@912_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@911 N_OUT9_Mn9@911_d N_OUT8_Mn9@911_g N_VSS_Mn9@911_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@910 N_OUT9_Mn9@910_d N_OUT8_Mn9@910_g N_VSS_Mn9@910_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@911 N_OUT9_Mp9@911_d N_OUT8_Mp9@911_g N_VDD_Mp9@911_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@910 N_OUT9_Mp9@910_d N_OUT8_Mp9@910_g N_VDD_Mp9@910_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@909 N_OUT9_Mn9@909_d N_OUT8_Mn9@909_g N_VSS_Mn9@909_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@908 N_OUT9_Mn9@908_d N_OUT8_Mn9@908_g N_VSS_Mn9@908_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@909 N_OUT9_Mp9@909_d N_OUT8_Mp9@909_g N_VDD_Mp9@909_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@908 N_OUT9_Mp9@908_d N_OUT8_Mp9@908_g N_VDD_Mp9@908_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@907 N_OUT9_Mn9@907_d N_OUT8_Mn9@907_g N_VSS_Mn9@907_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@906 N_OUT9_Mn9@906_d N_OUT8_Mn9@906_g N_VSS_Mn9@906_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@907 N_OUT9_Mp9@907_d N_OUT8_Mp9@907_g N_VDD_Mp9@907_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@906 N_OUT9_Mp9@906_d N_OUT8_Mp9@906_g N_VDD_Mp9@906_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@905 N_OUT9_Mn9@905_d N_OUT8_Mn9@905_g N_VSS_Mn9@905_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@904 N_OUT9_Mn9@904_d N_OUT8_Mn9@904_g N_VSS_Mn9@904_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@905 N_OUT9_Mp9@905_d N_OUT8_Mp9@905_g N_VDD_Mp9@905_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@904 N_OUT9_Mp9@904_d N_OUT8_Mp9@904_g N_VDD_Mp9@904_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@903 N_OUT9_Mn9@903_d N_OUT8_Mn9@903_g N_VSS_Mn9@903_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@902 N_OUT9_Mn9@902_d N_OUT8_Mn9@902_g N_VSS_Mn9@902_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@903 N_OUT9_Mp9@903_d N_OUT8_Mp9@903_g N_VDD_Mp9@903_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@902 N_OUT9_Mp9@902_d N_OUT8_Mp9@902_g N_VDD_Mp9@902_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@901 N_OUT9_Mn9@901_d N_OUT8_Mn9@901_g N_VSS_Mn9@901_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@900 N_OUT9_Mn9@900_d N_OUT8_Mn9@900_g N_VSS_Mn9@900_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@901 N_OUT9_Mp9@901_d N_OUT8_Mp9@901_g N_VDD_Mp9@901_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@900 N_OUT9_Mp9@900_d N_OUT8_Mp9@900_g N_VDD_Mp9@900_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@899 N_OUT9_Mn9@899_d N_OUT8_Mn9@899_g N_VSS_Mn9@899_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@898 N_OUT9_Mn9@898_d N_OUT8_Mn9@898_g N_VSS_Mn9@898_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@899 N_OUT9_Mp9@899_d N_OUT8_Mp9@899_g N_VDD_Mp9@899_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@898 N_OUT9_Mp9@898_d N_OUT8_Mp9@898_g N_VDD_Mp9@898_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@897 N_OUT9_Mn9@897_d N_OUT8_Mn9@897_g N_VSS_Mn9@897_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@896 N_OUT9_Mn9@896_d N_OUT8_Mn9@896_g N_VSS_Mn9@896_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@897 N_OUT9_Mp9@897_d N_OUT8_Mp9@897_g N_VDD_Mp9@897_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@896 N_OUT9_Mp9@896_d N_OUT8_Mp9@896_g N_VDD_Mp9@896_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@895 N_OUT9_Mn9@895_d N_OUT8_Mn9@895_g N_VSS_Mn9@895_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@894 N_OUT9_Mn9@894_d N_OUT8_Mn9@894_g N_VSS_Mn9@894_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@895 N_OUT9_Mp9@895_d N_OUT8_Mp9@895_g N_VDD_Mp9@895_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@894 N_OUT9_Mp9@894_d N_OUT8_Mp9@894_g N_VDD_Mp9@894_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@893 N_OUT9_Mn9@893_d N_OUT8_Mn9@893_g N_VSS_Mn9@893_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@892 N_OUT9_Mn9@892_d N_OUT8_Mn9@892_g N_VSS_Mn9@892_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@893 N_OUT9_Mp9@893_d N_OUT8_Mp9@893_g N_VDD_Mp9@893_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@892 N_OUT9_Mp9@892_d N_OUT8_Mp9@892_g N_VDD_Mp9@892_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@891 N_OUT9_Mn9@891_d N_OUT8_Mn9@891_g N_VSS_Mn9@891_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@890 N_OUT9_Mn9@890_d N_OUT8_Mn9@890_g N_VSS_Mn9@890_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@891 N_OUT9_Mp9@891_d N_OUT8_Mp9@891_g N_VDD_Mp9@891_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@890 N_OUT9_Mp9@890_d N_OUT8_Mp9@890_g N_VDD_Mp9@890_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@889 N_OUT9_Mn9@889_d N_OUT8_Mn9@889_g N_VSS_Mn9@889_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@888 N_OUT9_Mn9@888_d N_OUT8_Mn9@888_g N_VSS_Mn9@888_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@889 N_OUT9_Mp9@889_d N_OUT8_Mp9@889_g N_VDD_Mp9@889_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@888 N_OUT9_Mp9@888_d N_OUT8_Mp9@888_g N_VDD_Mp9@888_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@887 N_OUT9_Mn9@887_d N_OUT8_Mn9@887_g N_VSS_Mn9@887_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@886 N_OUT9_Mn9@886_d N_OUT8_Mn9@886_g N_VSS_Mn9@886_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@887 N_OUT9_Mp9@887_d N_OUT8_Mp9@887_g N_VDD_Mp9@887_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@886 N_OUT9_Mp9@886_d N_OUT8_Mp9@886_g N_VDD_Mp9@886_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@885 N_OUT9_Mn9@885_d N_OUT8_Mn9@885_g N_VSS_Mn9@885_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@884 N_OUT9_Mn9@884_d N_OUT8_Mn9@884_g N_VSS_Mn9@884_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@885 N_OUT9_Mp9@885_d N_OUT8_Mp9@885_g N_VDD_Mp9@885_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@884 N_OUT9_Mp9@884_d N_OUT8_Mp9@884_g N_VDD_Mp9@884_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@883 N_OUT9_Mn9@883_d N_OUT8_Mn9@883_g N_VSS_Mn9@883_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@882 N_OUT9_Mn9@882_d N_OUT8_Mn9@882_g N_VSS_Mn9@882_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@883 N_OUT9_Mp9@883_d N_OUT8_Mp9@883_g N_VDD_Mp9@883_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@882 N_OUT9_Mp9@882_d N_OUT8_Mp9@882_g N_VDD_Mp9@882_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@881 N_OUT9_Mn9@881_d N_OUT8_Mn9@881_g N_VSS_Mn9@881_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@880 N_OUT9_Mn9@880_d N_OUT8_Mn9@880_g N_VSS_Mn9@880_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@881 N_OUT9_Mp9@881_d N_OUT8_Mp9@881_g N_VDD_Mp9@881_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@880 N_OUT9_Mp9@880_d N_OUT8_Mp9@880_g N_VDD_Mp9@880_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@879 N_OUT9_Mn9@879_d N_OUT8_Mn9@879_g N_VSS_Mn9@879_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@878 N_OUT9_Mn9@878_d N_OUT8_Mn9@878_g N_VSS_Mn9@878_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@879 N_OUT9_Mp9@879_d N_OUT8_Mp9@879_g N_VDD_Mp9@879_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@878 N_OUT9_Mp9@878_d N_OUT8_Mp9@878_g N_VDD_Mp9@878_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@877 N_OUT9_Mn9@877_d N_OUT8_Mn9@877_g N_VSS_Mn9@877_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@876 N_OUT9_Mn9@876_d N_OUT8_Mn9@876_g N_VSS_Mn9@876_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@877 N_OUT9_Mp9@877_d N_OUT8_Mp9@877_g N_VDD_Mp9@877_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@876 N_OUT9_Mp9@876_d N_OUT8_Mp9@876_g N_VDD_Mp9@876_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@875 N_OUT9_Mn9@875_d N_OUT8_Mn9@875_g N_VSS_Mn9@875_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@874 N_OUT9_Mn9@874_d N_OUT8_Mn9@874_g N_VSS_Mn9@874_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@875 N_OUT9_Mp9@875_d N_OUT8_Mp9@875_g N_VDD_Mp9@875_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@874 N_OUT9_Mp9@874_d N_OUT8_Mp9@874_g N_VDD_Mp9@874_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@873 N_OUT9_Mn9@873_d N_OUT8_Mn9@873_g N_VSS_Mn9@873_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@872 N_OUT9_Mn9@872_d N_OUT8_Mn9@872_g N_VSS_Mn9@872_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@873 N_OUT9_Mp9@873_d N_OUT8_Mp9@873_g N_VDD_Mp9@873_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@872 N_OUT9_Mp9@872_d N_OUT8_Mp9@872_g N_VDD_Mp9@872_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@871 N_OUT9_Mn9@871_d N_OUT8_Mn9@871_g N_VSS_Mn9@871_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@870 N_OUT9_Mn9@870_d N_OUT8_Mn9@870_g N_VSS_Mn9@870_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@871 N_OUT9_Mp9@871_d N_OUT8_Mp9@871_g N_VDD_Mp9@871_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@870 N_OUT9_Mp9@870_d N_OUT8_Mp9@870_g N_VDD_Mp9@870_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@869 N_OUT9_Mn9@869_d N_OUT8_Mn9@869_g N_VSS_Mn9@869_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@868 N_OUT9_Mn9@868_d N_OUT8_Mn9@868_g N_VSS_Mn9@868_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@869 N_OUT9_Mp9@869_d N_OUT8_Mp9@869_g N_VDD_Mp9@869_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@868 N_OUT9_Mp9@868_d N_OUT8_Mp9@868_g N_VDD_Mp9@868_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@867 N_OUT9_Mn9@867_d N_OUT8_Mn9@867_g N_VSS_Mn9@867_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@866 N_OUT9_Mn9@866_d N_OUT8_Mn9@866_g N_VSS_Mn9@866_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@867 N_OUT9_Mp9@867_d N_OUT8_Mp9@867_g N_VDD_Mp9@867_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@866 N_OUT9_Mp9@866_d N_OUT8_Mp9@866_g N_VDD_Mp9@866_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@865 N_OUT9_Mn9@865_d N_OUT8_Mn9@865_g N_VSS_Mn9@865_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@864 N_OUT9_Mn9@864_d N_OUT8_Mn9@864_g N_VSS_Mn9@864_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@865 N_OUT9_Mp9@865_d N_OUT8_Mp9@865_g N_VDD_Mp9@865_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@864 N_OUT9_Mp9@864_d N_OUT8_Mp9@864_g N_VDD_Mp9@864_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@863 N_OUT9_Mn9@863_d N_OUT8_Mn9@863_g N_VSS_Mn9@863_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@862 N_OUT9_Mn9@862_d N_OUT8_Mn9@862_g N_VSS_Mn9@862_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@863 N_OUT9_Mp9@863_d N_OUT8_Mp9@863_g N_VDD_Mp9@863_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@862 N_OUT9_Mp9@862_d N_OUT8_Mp9@862_g N_VDD_Mp9@862_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@861 N_OUT9_Mn9@861_d N_OUT8_Mn9@861_g N_VSS_Mn9@861_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@860 N_OUT9_Mn9@860_d N_OUT8_Mn9@860_g N_VSS_Mn9@860_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@861 N_OUT9_Mp9@861_d N_OUT8_Mp9@861_g N_VDD_Mp9@861_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@860 N_OUT9_Mp9@860_d N_OUT8_Mp9@860_g N_VDD_Mp9@860_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@859 N_OUT9_Mn9@859_d N_OUT8_Mn9@859_g N_VSS_Mn9@859_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@858 N_OUT9_Mn9@858_d N_OUT8_Mn9@858_g N_VSS_Mn9@858_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@859 N_OUT9_Mp9@859_d N_OUT8_Mp9@859_g N_VDD_Mp9@859_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@858 N_OUT9_Mp9@858_d N_OUT8_Mp9@858_g N_VDD_Mp9@858_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@857 N_OUT9_Mn9@857_d N_OUT8_Mn9@857_g N_VSS_Mn9@857_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@856 N_OUT9_Mn9@856_d N_OUT8_Mn9@856_g N_VSS_Mn9@856_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@857 N_OUT9_Mp9@857_d N_OUT8_Mp9@857_g N_VDD_Mp9@857_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@856 N_OUT9_Mp9@856_d N_OUT8_Mp9@856_g N_VDD_Mp9@856_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@855 N_OUT9_Mn9@855_d N_OUT8_Mn9@855_g N_VSS_Mn9@855_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@854 N_OUT9_Mn9@854_d N_OUT8_Mn9@854_g N_VSS_Mn9@854_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@855 N_OUT9_Mp9@855_d N_OUT8_Mp9@855_g N_VDD_Mp9@855_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@854 N_OUT9_Mp9@854_d N_OUT8_Mp9@854_g N_VDD_Mp9@854_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@853 N_OUT9_Mn9@853_d N_OUT8_Mn9@853_g N_VSS_Mn9@853_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@852 N_OUT9_Mn9@852_d N_OUT8_Mn9@852_g N_VSS_Mn9@852_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@853 N_OUT9_Mp9@853_d N_OUT8_Mp9@853_g N_VDD_Mp9@853_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@852 N_OUT9_Mp9@852_d N_OUT8_Mp9@852_g N_VDD_Mp9@852_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@851 N_OUT9_Mn9@851_d N_OUT8_Mn9@851_g N_VSS_Mn9@851_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@850 N_OUT9_Mn9@850_d N_OUT8_Mn9@850_g N_VSS_Mn9@850_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@851 N_OUT9_Mp9@851_d N_OUT8_Mp9@851_g N_VDD_Mp9@851_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@850 N_OUT9_Mp9@850_d N_OUT8_Mp9@850_g N_VDD_Mp9@850_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@849 N_OUT9_Mn9@849_d N_OUT8_Mn9@849_g N_VSS_Mn9@849_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@848 N_OUT9_Mn9@848_d N_OUT8_Mn9@848_g N_VSS_Mn9@848_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@849 N_OUT9_Mp9@849_d N_OUT8_Mp9@849_g N_VDD_Mp9@849_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@848 N_OUT9_Mp9@848_d N_OUT8_Mp9@848_g N_VDD_Mp9@848_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@847 N_OUT9_Mn9@847_d N_OUT8_Mn9@847_g N_VSS_Mn9@847_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@846 N_OUT9_Mn9@846_d N_OUT8_Mn9@846_g N_VSS_Mn9@846_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@847 N_OUT9_Mp9@847_d N_OUT8_Mp9@847_g N_VDD_Mp9@847_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@846 N_OUT9_Mp9@846_d N_OUT8_Mp9@846_g N_VDD_Mp9@846_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@845 N_OUT9_Mn9@845_d N_OUT8_Mn9@845_g N_VSS_Mn9@845_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@844 N_OUT9_Mn9@844_d N_OUT8_Mn9@844_g N_VSS_Mn9@844_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@845 N_OUT9_Mp9@845_d N_OUT8_Mp9@845_g N_VDD_Mp9@845_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@844 N_OUT9_Mp9@844_d N_OUT8_Mp9@844_g N_VDD_Mp9@844_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@843 N_OUT9_Mn9@843_d N_OUT8_Mn9@843_g N_VSS_Mn9@843_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@842 N_OUT9_Mn9@842_d N_OUT8_Mn9@842_g N_VSS_Mn9@842_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@843 N_OUT9_Mp9@843_d N_OUT8_Mp9@843_g N_VDD_Mp9@843_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@842 N_OUT9_Mp9@842_d N_OUT8_Mp9@842_g N_VDD_Mp9@842_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@841 N_OUT9_Mn9@841_d N_OUT8_Mn9@841_g N_VSS_Mn9@841_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@840 N_OUT9_Mn9@840_d N_OUT8_Mn9@840_g N_VSS_Mn9@840_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@841 N_OUT9_Mp9@841_d N_OUT8_Mp9@841_g N_VDD_Mp9@841_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@840 N_OUT9_Mp9@840_d N_OUT8_Mp9@840_g N_VDD_Mp9@840_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@839 N_OUT9_Mn9@839_d N_OUT8_Mn9@839_g N_VSS_Mn9@839_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@838 N_OUT9_Mn9@838_d N_OUT8_Mn9@838_g N_VSS_Mn9@838_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@839 N_OUT9_Mp9@839_d N_OUT8_Mp9@839_g N_VDD_Mp9@839_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@838 N_OUT9_Mp9@838_d N_OUT8_Mp9@838_g N_VDD_Mp9@838_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@837 N_OUT9_Mn9@837_d N_OUT8_Mn9@837_g N_VSS_Mn9@837_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@836 N_OUT9_Mn9@836_d N_OUT8_Mn9@836_g N_VSS_Mn9@836_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@837 N_OUT9_Mp9@837_d N_OUT8_Mp9@837_g N_VDD_Mp9@837_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@836 N_OUT9_Mp9@836_d N_OUT8_Mp9@836_g N_VDD_Mp9@836_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@835 N_OUT9_Mn9@835_d N_OUT8_Mn9@835_g N_VSS_Mn9@835_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@834 N_OUT9_Mn9@834_d N_OUT8_Mn9@834_g N_VSS_Mn9@834_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@835 N_OUT9_Mp9@835_d N_OUT8_Mp9@835_g N_VDD_Mp9@835_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@834 N_OUT9_Mp9@834_d N_OUT8_Mp9@834_g N_VDD_Mp9@834_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@833 N_OUT9_Mn9@833_d N_OUT8_Mn9@833_g N_VSS_Mn9@833_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@832 N_OUT9_Mn9@832_d N_OUT8_Mn9@832_g N_VSS_Mn9@832_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@833 N_OUT9_Mp9@833_d N_OUT8_Mp9@833_g N_VDD_Mp9@833_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@832 N_OUT9_Mp9@832_d N_OUT8_Mp9@832_g N_VDD_Mp9@832_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@831 N_OUT9_Mn9@831_d N_OUT8_Mn9@831_g N_VSS_Mn9@831_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@830 N_OUT9_Mn9@830_d N_OUT8_Mn9@830_g N_VSS_Mn9@830_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@831 N_OUT9_Mp9@831_d N_OUT8_Mp9@831_g N_VDD_Mp9@831_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@830 N_OUT9_Mp9@830_d N_OUT8_Mp9@830_g N_VDD_Mp9@830_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@829 N_OUT9_Mn9@829_d N_OUT8_Mn9@829_g N_VSS_Mn9@829_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@828 N_OUT9_Mn9@828_d N_OUT8_Mn9@828_g N_VSS_Mn9@828_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@829 N_OUT9_Mp9@829_d N_OUT8_Mp9@829_g N_VDD_Mp9@829_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@828 N_OUT9_Mp9@828_d N_OUT8_Mp9@828_g N_VDD_Mp9@828_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@827 N_OUT9_Mn9@827_d N_OUT8_Mn9@827_g N_VSS_Mn9@827_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@826 N_OUT9_Mn9@826_d N_OUT8_Mn9@826_g N_VSS_Mn9@826_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@827 N_OUT9_Mp9@827_d N_OUT8_Mp9@827_g N_VDD_Mp9@827_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@826 N_OUT9_Mp9@826_d N_OUT8_Mp9@826_g N_VDD_Mp9@826_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@825 N_OUT9_Mn9@825_d N_OUT8_Mn9@825_g N_VSS_Mn9@825_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@824 N_OUT9_Mn9@824_d N_OUT8_Mn9@824_g N_VSS_Mn9@824_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@825 N_OUT9_Mp9@825_d N_OUT8_Mp9@825_g N_VDD_Mp9@825_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@824 N_OUT9_Mp9@824_d N_OUT8_Mp9@824_g N_VDD_Mp9@824_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@823 N_OUT9_Mn9@823_d N_OUT8_Mn9@823_g N_VSS_Mn9@823_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@822 N_OUT9_Mn9@822_d N_OUT8_Mn9@822_g N_VSS_Mn9@822_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@823 N_OUT9_Mp9@823_d N_OUT8_Mp9@823_g N_VDD_Mp9@823_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@822 N_OUT9_Mp9@822_d N_OUT8_Mp9@822_g N_VDD_Mp9@822_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@821 N_OUT9_Mn9@821_d N_OUT8_Mn9@821_g N_VSS_Mn9@821_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@820 N_OUT9_Mn9@820_d N_OUT8_Mn9@820_g N_VSS_Mn9@820_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@821 N_OUT9_Mp9@821_d N_OUT8_Mp9@821_g N_VDD_Mp9@821_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@820 N_OUT9_Mp9@820_d N_OUT8_Mp9@820_g N_VDD_Mp9@820_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@819 N_OUT9_Mn9@819_d N_OUT8_Mn9@819_g N_VSS_Mn9@819_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@818 N_OUT9_Mn9@818_d N_OUT8_Mn9@818_g N_VSS_Mn9@818_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@819 N_OUT9_Mp9@819_d N_OUT8_Mp9@819_g N_VDD_Mp9@819_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@818 N_OUT9_Mp9@818_d N_OUT8_Mp9@818_g N_VDD_Mp9@818_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@817 N_OUT9_Mn9@817_d N_OUT8_Mn9@817_g N_VSS_Mn9@817_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@816 N_OUT9_Mn9@816_d N_OUT8_Mn9@816_g N_VSS_Mn9@816_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@817 N_OUT9_Mp9@817_d N_OUT8_Mp9@817_g N_VDD_Mp9@817_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@816 N_OUT9_Mp9@816_d N_OUT8_Mp9@816_g N_VDD_Mp9@816_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@815 N_OUT9_Mn9@815_d N_OUT8_Mn9@815_g N_VSS_Mn9@815_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@814 N_OUT9_Mn9@814_d N_OUT8_Mn9@814_g N_VSS_Mn9@814_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@815 N_OUT9_Mp9@815_d N_OUT8_Mp9@815_g N_VDD_Mp9@815_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@814 N_OUT9_Mp9@814_d N_OUT8_Mp9@814_g N_VDD_Mp9@814_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@813 N_OUT9_Mn9@813_d N_OUT8_Mn9@813_g N_VSS_Mn9@813_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@812 N_OUT9_Mn9@812_d N_OUT8_Mn9@812_g N_VSS_Mn9@812_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@813 N_OUT9_Mp9@813_d N_OUT8_Mp9@813_g N_VDD_Mp9@813_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@812 N_OUT9_Mp9@812_d N_OUT8_Mp9@812_g N_VDD_Mp9@812_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@811 N_OUT9_Mn9@811_d N_OUT8_Mn9@811_g N_VSS_Mn9@811_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@810 N_OUT9_Mn9@810_d N_OUT8_Mn9@810_g N_VSS_Mn9@810_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@811 N_OUT9_Mp9@811_d N_OUT8_Mp9@811_g N_VDD_Mp9@811_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@810 N_OUT9_Mp9@810_d N_OUT8_Mp9@810_g N_VDD_Mp9@810_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@809 N_OUT9_Mn9@809_d N_OUT8_Mn9@809_g N_VSS_Mn9@809_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@808 N_OUT9_Mn9@808_d N_OUT8_Mn9@808_g N_VSS_Mn9@808_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@809 N_OUT9_Mp9@809_d N_OUT8_Mp9@809_g N_VDD_Mp9@809_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@808 N_OUT9_Mp9@808_d N_OUT8_Mp9@808_g N_VDD_Mp9@808_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@807 N_OUT9_Mn9@807_d N_OUT8_Mn9@807_g N_VSS_Mn9@807_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@806 N_OUT9_Mn9@806_d N_OUT8_Mn9@806_g N_VSS_Mn9@806_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@807 N_OUT9_Mp9@807_d N_OUT8_Mp9@807_g N_VDD_Mp9@807_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@806 N_OUT9_Mp9@806_d N_OUT8_Mp9@806_g N_VDD_Mp9@806_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@805 N_OUT9_Mn9@805_d N_OUT8_Mn9@805_g N_VSS_Mn9@805_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@804 N_OUT9_Mn9@804_d N_OUT8_Mn9@804_g N_VSS_Mn9@804_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@805 N_OUT9_Mp9@805_d N_OUT8_Mp9@805_g N_VDD_Mp9@805_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@804 N_OUT9_Mp9@804_d N_OUT8_Mp9@804_g N_VDD_Mp9@804_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@803 N_OUT9_Mn9@803_d N_OUT8_Mn9@803_g N_VSS_Mn9@803_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@802 N_OUT9_Mn9@802_d N_OUT8_Mn9@802_g N_VSS_Mn9@802_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@803 N_OUT9_Mp9@803_d N_OUT8_Mp9@803_g N_VDD_Mp9@803_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@802 N_OUT9_Mp9@802_d N_OUT8_Mp9@802_g N_VDD_Mp9@802_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@801 N_OUT9_Mn9@801_d N_OUT8_Mn9@801_g N_VSS_Mn9@801_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@800 N_OUT9_Mn9@800_d N_OUT8_Mn9@800_g N_VSS_Mn9@800_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@801 N_OUT9_Mp9@801_d N_OUT8_Mp9@801_g N_VDD_Mp9@801_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@800 N_OUT9_Mp9@800_d N_OUT8_Mp9@800_g N_VDD_Mp9@800_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@799 N_OUT9_Mn9@799_d N_OUT8_Mn9@799_g N_VSS_Mn9@799_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@798 N_OUT9_Mn9@798_d N_OUT8_Mn9@798_g N_VSS_Mn9@798_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@799 N_OUT9_Mp9@799_d N_OUT8_Mp9@799_g N_VDD_Mp9@799_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@798 N_OUT9_Mp9@798_d N_OUT8_Mp9@798_g N_VDD_Mp9@798_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@797 N_OUT9_Mn9@797_d N_OUT8_Mn9@797_g N_VSS_Mn9@797_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@796 N_OUT9_Mn9@796_d N_OUT8_Mn9@796_g N_VSS_Mn9@796_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@797 N_OUT9_Mp9@797_d N_OUT8_Mp9@797_g N_VDD_Mp9@797_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@796 N_OUT9_Mp9@796_d N_OUT8_Mp9@796_g N_VDD_Mp9@796_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@795 N_OUT9_Mn9@795_d N_OUT8_Mn9@795_g N_VSS_Mn9@795_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@794 N_OUT9_Mn9@794_d N_OUT8_Mn9@794_g N_VSS_Mn9@794_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@795 N_OUT9_Mp9@795_d N_OUT8_Mp9@795_g N_VDD_Mp9@795_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@794 N_OUT9_Mp9@794_d N_OUT8_Mp9@794_g N_VDD_Mp9@794_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@793 N_OUT9_Mn9@793_d N_OUT8_Mn9@793_g N_VSS_Mn9@793_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@792 N_OUT9_Mn9@792_d N_OUT8_Mn9@792_g N_VSS_Mn9@792_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@793 N_OUT9_Mp9@793_d N_OUT8_Mp9@793_g N_VDD_Mp9@793_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@792 N_OUT9_Mp9@792_d N_OUT8_Mp9@792_g N_VDD_Mp9@792_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@791 N_OUT9_Mn9@791_d N_OUT8_Mn9@791_g N_VSS_Mn9@791_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@790 N_OUT9_Mn9@790_d N_OUT8_Mn9@790_g N_VSS_Mn9@790_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@791 N_OUT9_Mp9@791_d N_OUT8_Mp9@791_g N_VDD_Mp9@791_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@790 N_OUT9_Mp9@790_d N_OUT8_Mp9@790_g N_VDD_Mp9@790_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@789 N_OUT9_Mn9@789_d N_OUT8_Mn9@789_g N_VSS_Mn9@789_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@788 N_OUT9_Mn9@788_d N_OUT8_Mn9@788_g N_VSS_Mn9@788_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@789 N_OUT9_Mp9@789_d N_OUT8_Mp9@789_g N_VDD_Mp9@789_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@788 N_OUT9_Mp9@788_d N_OUT8_Mp9@788_g N_VDD_Mp9@788_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@787 N_OUT9_Mn9@787_d N_OUT8_Mn9@787_g N_VSS_Mn9@787_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@786 N_OUT9_Mn9@786_d N_OUT8_Mn9@786_g N_VSS_Mn9@786_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@787 N_OUT9_Mp9@787_d N_OUT8_Mp9@787_g N_VDD_Mp9@787_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@786 N_OUT9_Mp9@786_d N_OUT8_Mp9@786_g N_VDD_Mp9@786_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@785 N_OUT9_Mn9@785_d N_OUT8_Mn9@785_g N_VSS_Mn9@785_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@784 N_OUT9_Mn9@784_d N_OUT8_Mn9@784_g N_VSS_Mn9@784_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@785 N_OUT9_Mp9@785_d N_OUT8_Mp9@785_g N_VDD_Mp9@785_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@784 N_OUT9_Mp9@784_d N_OUT8_Mp9@784_g N_VDD_Mp9@784_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@783 N_OUT9_Mn9@783_d N_OUT8_Mn9@783_g N_VSS_Mn9@783_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@782 N_OUT9_Mn9@782_d N_OUT8_Mn9@782_g N_VSS_Mn9@782_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@783 N_OUT9_Mp9@783_d N_OUT8_Mp9@783_g N_VDD_Mp9@783_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@782 N_OUT9_Mp9@782_d N_OUT8_Mp9@782_g N_VDD_Mp9@782_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@781 N_OUT9_Mn9@781_d N_OUT8_Mn9@781_g N_VSS_Mn9@781_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@780 N_OUT9_Mn9@780_d N_OUT8_Mn9@780_g N_VSS_Mn9@780_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@781 N_OUT9_Mp9@781_d N_OUT8_Mp9@781_g N_VDD_Mp9@781_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@780 N_OUT9_Mp9@780_d N_OUT8_Mp9@780_g N_VDD_Mp9@780_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@779 N_OUT9_Mn9@779_d N_OUT8_Mn9@779_g N_VSS_Mn9@779_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@778 N_OUT9_Mn9@778_d N_OUT8_Mn9@778_g N_VSS_Mn9@778_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@779 N_OUT9_Mp9@779_d N_OUT8_Mp9@779_g N_VDD_Mp9@779_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@778 N_OUT9_Mp9@778_d N_OUT8_Mp9@778_g N_VDD_Mp9@778_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@777 N_OUT9_Mn9@777_d N_OUT8_Mn9@777_g N_VSS_Mn9@777_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@776 N_OUT9_Mn9@776_d N_OUT8_Mn9@776_g N_VSS_Mn9@776_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@777 N_OUT9_Mp9@777_d N_OUT8_Mp9@777_g N_VDD_Mp9@777_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@776 N_OUT9_Mp9@776_d N_OUT8_Mp9@776_g N_VDD_Mp9@776_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@775 N_OUT9_Mn9@775_d N_OUT8_Mn9@775_g N_VSS_Mn9@775_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@774 N_OUT9_Mn9@774_d N_OUT8_Mn9@774_g N_VSS_Mn9@774_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@775 N_OUT9_Mp9@775_d N_OUT8_Mp9@775_g N_VDD_Mp9@775_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@774 N_OUT9_Mp9@774_d N_OUT8_Mp9@774_g N_VDD_Mp9@774_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@773 N_OUT9_Mn9@773_d N_OUT8_Mn9@773_g N_VSS_Mn9@773_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@772 N_OUT9_Mn9@772_d N_OUT8_Mn9@772_g N_VSS_Mn9@772_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@773 N_OUT9_Mp9@773_d N_OUT8_Mp9@773_g N_VDD_Mp9@773_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@772 N_OUT9_Mp9@772_d N_OUT8_Mp9@772_g N_VDD_Mp9@772_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@771 N_OUT9_Mn9@771_d N_OUT8_Mn9@771_g N_VSS_Mn9@771_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@770 N_OUT9_Mn9@770_d N_OUT8_Mn9@770_g N_VSS_Mn9@770_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@771 N_OUT9_Mp9@771_d N_OUT8_Mp9@771_g N_VDD_Mp9@771_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@770 N_OUT9_Mp9@770_d N_OUT8_Mp9@770_g N_VDD_Mp9@770_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@769 N_OUT9_Mn9@769_d N_OUT8_Mn9@769_g N_VSS_Mn9@769_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@768 N_OUT9_Mn9@768_d N_OUT8_Mn9@768_g N_VSS_Mn9@768_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@769 N_OUT9_Mp9@769_d N_OUT8_Mp9@769_g N_VDD_Mp9@769_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@768 N_OUT9_Mp9@768_d N_OUT8_Mp9@768_g N_VDD_Mp9@768_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@767 N_OUT9_Mn9@767_d N_OUT8_Mn9@767_g N_VSS_Mn9@767_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@766 N_OUT9_Mn9@766_d N_OUT8_Mn9@766_g N_VSS_Mn9@766_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@767 N_OUT9_Mp9@767_d N_OUT8_Mp9@767_g N_VDD_Mp9@767_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@766 N_OUT9_Mp9@766_d N_OUT8_Mp9@766_g N_VDD_Mp9@766_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@765 N_OUT9_Mn9@765_d N_OUT8_Mn9@765_g N_VSS_Mn9@765_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@764 N_OUT9_Mn9@764_d N_OUT8_Mn9@764_g N_VSS_Mn9@764_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@765 N_OUT9_Mp9@765_d N_OUT8_Mp9@765_g N_VDD_Mp9@765_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@764 N_OUT9_Mp9@764_d N_OUT8_Mp9@764_g N_VDD_Mp9@764_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@763 N_OUT9_Mn9@763_d N_OUT8_Mn9@763_g N_VSS_Mn9@763_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@762 N_OUT9_Mn9@762_d N_OUT8_Mn9@762_g N_VSS_Mn9@762_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@763 N_OUT9_Mp9@763_d N_OUT8_Mp9@763_g N_VDD_Mp9@763_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@762 N_OUT9_Mp9@762_d N_OUT8_Mp9@762_g N_VDD_Mp9@762_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@761 N_OUT9_Mn9@761_d N_OUT8_Mn9@761_g N_VSS_Mn9@761_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@760 N_OUT9_Mn9@760_d N_OUT8_Mn9@760_g N_VSS_Mn9@760_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@761 N_OUT9_Mp9@761_d N_OUT8_Mp9@761_g N_VDD_Mp9@761_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@760 N_OUT9_Mp9@760_d N_OUT8_Mp9@760_g N_VDD_Mp9@760_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@759 N_OUT9_Mn9@759_d N_OUT8_Mn9@759_g N_VSS_Mn9@759_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@758 N_OUT9_Mn9@758_d N_OUT8_Mn9@758_g N_VSS_Mn9@758_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@759 N_OUT9_Mp9@759_d N_OUT8_Mp9@759_g N_VDD_Mp9@759_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@758 N_OUT9_Mp9@758_d N_OUT8_Mp9@758_g N_VDD_Mp9@758_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@757 N_OUT9_Mn9@757_d N_OUT8_Mn9@757_g N_VSS_Mn9@757_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@756 N_OUT9_Mn9@756_d N_OUT8_Mn9@756_g N_VSS_Mn9@756_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@757 N_OUT9_Mp9@757_d N_OUT8_Mp9@757_g N_VDD_Mp9@757_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@756 N_OUT9_Mp9@756_d N_OUT8_Mp9@756_g N_VDD_Mp9@756_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@755 N_OUT9_Mn9@755_d N_OUT8_Mn9@755_g N_VSS_Mn9@755_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@754 N_OUT9_Mn9@754_d N_OUT8_Mn9@754_g N_VSS_Mn9@754_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@755 N_OUT9_Mp9@755_d N_OUT8_Mp9@755_g N_VDD_Mp9@755_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@754 N_OUT9_Mp9@754_d N_OUT8_Mp9@754_g N_VDD_Mp9@754_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@753 N_OUT9_Mn9@753_d N_OUT8_Mn9@753_g N_VSS_Mn9@753_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@752 N_OUT9_Mn9@752_d N_OUT8_Mn9@752_g N_VSS_Mn9@752_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@753 N_OUT9_Mp9@753_d N_OUT8_Mp9@753_g N_VDD_Mp9@753_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@752 N_OUT9_Mp9@752_d N_OUT8_Mp9@752_g N_VDD_Mp9@752_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@751 N_OUT9_Mn9@751_d N_OUT8_Mn9@751_g N_VSS_Mn9@751_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@750 N_OUT9_Mn9@750_d N_OUT8_Mn9@750_g N_VSS_Mn9@750_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@751 N_OUT9_Mp9@751_d N_OUT8_Mp9@751_g N_VDD_Mp9@751_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@750 N_OUT9_Mp9@750_d N_OUT8_Mp9@750_g N_VDD_Mp9@750_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@749 N_OUT9_Mn9@749_d N_OUT8_Mn9@749_g N_VSS_Mn9@749_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@748 N_OUT9_Mn9@748_d N_OUT8_Mn9@748_g N_VSS_Mn9@748_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@749 N_OUT9_Mp9@749_d N_OUT8_Mp9@749_g N_VDD_Mp9@749_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@748 N_OUT9_Mp9@748_d N_OUT8_Mp9@748_g N_VDD_Mp9@748_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@747 N_OUT9_Mn9@747_d N_OUT8_Mn9@747_g N_VSS_Mn9@747_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@746 N_OUT9_Mn9@746_d N_OUT8_Mn9@746_g N_VSS_Mn9@746_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@747 N_OUT9_Mp9@747_d N_OUT8_Mp9@747_g N_VDD_Mp9@747_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@746 N_OUT9_Mp9@746_d N_OUT8_Mp9@746_g N_VDD_Mp9@746_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@745 N_OUT9_Mn9@745_d N_OUT8_Mn9@745_g N_VSS_Mn9@745_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@744 N_OUT9_Mn9@744_d N_OUT8_Mn9@744_g N_VSS_Mn9@744_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@745 N_OUT9_Mp9@745_d N_OUT8_Mp9@745_g N_VDD_Mp9@745_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@744 N_OUT9_Mp9@744_d N_OUT8_Mp9@744_g N_VDD_Mp9@744_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@743 N_OUT9_Mn9@743_d N_OUT8_Mn9@743_g N_VSS_Mn9@743_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@742 N_OUT9_Mn9@742_d N_OUT8_Mn9@742_g N_VSS_Mn9@742_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@743 N_OUT9_Mp9@743_d N_OUT8_Mp9@743_g N_VDD_Mp9@743_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@742 N_OUT9_Mp9@742_d N_OUT8_Mp9@742_g N_VDD_Mp9@742_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@741 N_OUT9_Mn9@741_d N_OUT8_Mn9@741_g N_VSS_Mn9@741_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@740 N_OUT9_Mn9@740_d N_OUT8_Mn9@740_g N_VSS_Mn9@740_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@741 N_OUT9_Mp9@741_d N_OUT8_Mp9@741_g N_VDD_Mp9@741_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@740 N_OUT9_Mp9@740_d N_OUT8_Mp9@740_g N_VDD_Mp9@740_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@739 N_OUT9_Mn9@739_d N_OUT8_Mn9@739_g N_VSS_Mn9@739_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@738 N_OUT9_Mn9@738_d N_OUT8_Mn9@738_g N_VSS_Mn9@738_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@739 N_OUT9_Mp9@739_d N_OUT8_Mp9@739_g N_VDD_Mp9@739_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@738 N_OUT9_Mp9@738_d N_OUT8_Mp9@738_g N_VDD_Mp9@738_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@737 N_OUT9_Mn9@737_d N_OUT8_Mn9@737_g N_VSS_Mn9@737_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@736 N_OUT9_Mn9@736_d N_OUT8_Mn9@736_g N_VSS_Mn9@736_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@737 N_OUT9_Mp9@737_d N_OUT8_Mp9@737_g N_VDD_Mp9@737_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@736 N_OUT9_Mp9@736_d N_OUT8_Mp9@736_g N_VDD_Mp9@736_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@735 N_OUT9_Mn9@735_d N_OUT8_Mn9@735_g N_VSS_Mn9@735_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@734 N_OUT9_Mn9@734_d N_OUT8_Mn9@734_g N_VSS_Mn9@734_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@735 N_OUT9_Mp9@735_d N_OUT8_Mp9@735_g N_VDD_Mp9@735_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@734 N_OUT9_Mp9@734_d N_OUT8_Mp9@734_g N_VDD_Mp9@734_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@733 N_OUT9_Mn9@733_d N_OUT8_Mn9@733_g N_VSS_Mn9@733_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@732 N_OUT9_Mn9@732_d N_OUT8_Mn9@732_g N_VSS_Mn9@732_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@733 N_OUT9_Mp9@733_d N_OUT8_Mp9@733_g N_VDD_Mp9@733_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@732 N_OUT9_Mp9@732_d N_OUT8_Mp9@732_g N_VDD_Mp9@732_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@731 N_OUT9_Mn9@731_d N_OUT8_Mn9@731_g N_VSS_Mn9@731_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@730 N_OUT9_Mn9@730_d N_OUT8_Mn9@730_g N_VSS_Mn9@730_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@731 N_OUT9_Mp9@731_d N_OUT8_Mp9@731_g N_VDD_Mp9@731_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@730 N_OUT9_Mp9@730_d N_OUT8_Mp9@730_g N_VDD_Mp9@730_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@729 N_OUT9_Mn9@729_d N_OUT8_Mn9@729_g N_VSS_Mn9@729_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@728 N_OUT9_Mn9@728_d N_OUT8_Mn9@728_g N_VSS_Mn9@728_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@729 N_OUT9_Mp9@729_d N_OUT8_Mp9@729_g N_VDD_Mp9@729_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@728 N_OUT9_Mp9@728_d N_OUT8_Mp9@728_g N_VDD_Mp9@728_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@727 N_OUT9_Mn9@727_d N_OUT8_Mn9@727_g N_VSS_Mn9@727_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@726 N_OUT9_Mn9@726_d N_OUT8_Mn9@726_g N_VSS_Mn9@726_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@727 N_OUT9_Mp9@727_d N_OUT8_Mp9@727_g N_VDD_Mp9@727_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@726 N_OUT9_Mp9@726_d N_OUT8_Mp9@726_g N_VDD_Mp9@726_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@725 N_OUT9_Mn9@725_d N_OUT8_Mn9@725_g N_VSS_Mn9@725_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@724 N_OUT9_Mn9@724_d N_OUT8_Mn9@724_g N_VSS_Mn9@724_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@725 N_OUT9_Mp9@725_d N_OUT8_Mp9@725_g N_VDD_Mp9@725_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@724 N_OUT9_Mp9@724_d N_OUT8_Mp9@724_g N_VDD_Mp9@724_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@723 N_OUT9_Mn9@723_d N_OUT8_Mn9@723_g N_VSS_Mn9@723_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@722 N_OUT9_Mn9@722_d N_OUT8_Mn9@722_g N_VSS_Mn9@722_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@723 N_OUT9_Mp9@723_d N_OUT8_Mp9@723_g N_VDD_Mp9@723_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@722 N_OUT9_Mp9@722_d N_OUT8_Mp9@722_g N_VDD_Mp9@722_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@721 N_OUT9_Mn9@721_d N_OUT8_Mn9@721_g N_VSS_Mn9@721_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@720 N_OUT9_Mn9@720_d N_OUT8_Mn9@720_g N_VSS_Mn9@720_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@721 N_OUT9_Mp9@721_d N_OUT8_Mp9@721_g N_VDD_Mp9@721_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@720 N_OUT9_Mp9@720_d N_OUT8_Mp9@720_g N_VDD_Mp9@720_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@719 N_OUT9_Mn9@719_d N_OUT8_Mn9@719_g N_VSS_Mn9@719_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@718 N_OUT9_Mn9@718_d N_OUT8_Mn9@718_g N_VSS_Mn9@718_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@719 N_OUT9_Mp9@719_d N_OUT8_Mp9@719_g N_VDD_Mp9@719_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@718 N_OUT9_Mp9@718_d N_OUT8_Mp9@718_g N_VDD_Mp9@718_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@717 N_OUT9_Mn9@717_d N_OUT8_Mn9@717_g N_VSS_Mn9@717_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@716 N_OUT9_Mn9@716_d N_OUT8_Mn9@716_g N_VSS_Mn9@716_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@717 N_OUT9_Mp9@717_d N_OUT8_Mp9@717_g N_VDD_Mp9@717_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@716 N_OUT9_Mp9@716_d N_OUT8_Mp9@716_g N_VDD_Mp9@716_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@715 N_OUT9_Mn9@715_d N_OUT8_Mn9@715_g N_VSS_Mn9@715_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@714 N_OUT9_Mn9@714_d N_OUT8_Mn9@714_g N_VSS_Mn9@714_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@715 N_OUT9_Mp9@715_d N_OUT8_Mp9@715_g N_VDD_Mp9@715_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@714 N_OUT9_Mp9@714_d N_OUT8_Mp9@714_g N_VDD_Mp9@714_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@713 N_OUT9_Mn9@713_d N_OUT8_Mn9@713_g N_VSS_Mn9@713_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@712 N_OUT9_Mn9@712_d N_OUT8_Mn9@712_g N_VSS_Mn9@712_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@713 N_OUT9_Mp9@713_d N_OUT8_Mp9@713_g N_VDD_Mp9@713_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@712 N_OUT9_Mp9@712_d N_OUT8_Mp9@712_g N_VDD_Mp9@712_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@711 N_OUT9_Mn9@711_d N_OUT8_Mn9@711_g N_VSS_Mn9@711_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@710 N_OUT9_Mn9@710_d N_OUT8_Mn9@710_g N_VSS_Mn9@710_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@711 N_OUT9_Mp9@711_d N_OUT8_Mp9@711_g N_VDD_Mp9@711_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@710 N_OUT9_Mp9@710_d N_OUT8_Mp9@710_g N_VDD_Mp9@710_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@709 N_OUT9_Mn9@709_d N_OUT8_Mn9@709_g N_VSS_Mn9@709_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@708 N_OUT9_Mn9@708_d N_OUT8_Mn9@708_g N_VSS_Mn9@708_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@709 N_OUT9_Mp9@709_d N_OUT8_Mp9@709_g N_VDD_Mp9@709_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@708 N_OUT9_Mp9@708_d N_OUT8_Mp9@708_g N_VDD_Mp9@708_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@707 N_OUT9_Mn9@707_d N_OUT8_Mn9@707_g N_VSS_Mn9@707_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@706 N_OUT9_Mn9@706_d N_OUT8_Mn9@706_g N_VSS_Mn9@706_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@707 N_OUT9_Mp9@707_d N_OUT8_Mp9@707_g N_VDD_Mp9@707_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@706 N_OUT9_Mp9@706_d N_OUT8_Mp9@706_g N_VDD_Mp9@706_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@705 N_OUT9_Mn9@705_d N_OUT8_Mn9@705_g N_VSS_Mn9@705_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@704 N_OUT9_Mn9@704_d N_OUT8_Mn9@704_g N_VSS_Mn9@704_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@705 N_OUT9_Mp9@705_d N_OUT8_Mp9@705_g N_VDD_Mp9@705_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@704 N_OUT9_Mp9@704_d N_OUT8_Mp9@704_g N_VDD_Mp9@704_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@703 N_OUT9_Mn9@703_d N_OUT8_Mn9@703_g N_VSS_Mn9@703_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@702 N_OUT9_Mn9@702_d N_OUT8_Mn9@702_g N_VSS_Mn9@702_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@703 N_OUT9_Mp9@703_d N_OUT8_Mp9@703_g N_VDD_Mp9@703_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@702 N_OUT9_Mp9@702_d N_OUT8_Mp9@702_g N_VDD_Mp9@702_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@701 N_OUT9_Mn9@701_d N_OUT8_Mn9@701_g N_VSS_Mn9@701_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@700 N_OUT9_Mn9@700_d N_OUT8_Mn9@700_g N_VSS_Mn9@700_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@701 N_OUT9_Mp9@701_d N_OUT8_Mp9@701_g N_VDD_Mp9@701_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@700 N_OUT9_Mp9@700_d N_OUT8_Mp9@700_g N_VDD_Mp9@700_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@699 N_OUT9_Mn9@699_d N_OUT8_Mn9@699_g N_VSS_Mn9@699_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@698 N_OUT9_Mn9@698_d N_OUT8_Mn9@698_g N_VSS_Mn9@698_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@699 N_OUT9_Mp9@699_d N_OUT8_Mp9@699_g N_VDD_Mp9@699_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@698 N_OUT9_Mp9@698_d N_OUT8_Mp9@698_g N_VDD_Mp9@698_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@697 N_OUT9_Mn9@697_d N_OUT8_Mn9@697_g N_VSS_Mn9@697_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@696 N_OUT9_Mn9@696_d N_OUT8_Mn9@696_g N_VSS_Mn9@696_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@697 N_OUT9_Mp9@697_d N_OUT8_Mp9@697_g N_VDD_Mp9@697_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@696 N_OUT9_Mp9@696_d N_OUT8_Mp9@696_g N_VDD_Mp9@696_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@695 N_OUT9_Mn9@695_d N_OUT8_Mn9@695_g N_VSS_Mn9@695_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@694 N_OUT9_Mn9@694_d N_OUT8_Mn9@694_g N_VSS_Mn9@694_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@695 N_OUT9_Mp9@695_d N_OUT8_Mp9@695_g N_VDD_Mp9@695_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@694 N_OUT9_Mp9@694_d N_OUT8_Mp9@694_g N_VDD_Mp9@694_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@693 N_OUT9_Mn9@693_d N_OUT8_Mn9@693_g N_VSS_Mn9@693_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@692 N_OUT9_Mn9@692_d N_OUT8_Mn9@692_g N_VSS_Mn9@692_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@693 N_OUT9_Mp9@693_d N_OUT8_Mp9@693_g N_VDD_Mp9@693_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@692 N_OUT9_Mp9@692_d N_OUT8_Mp9@692_g N_VDD_Mp9@692_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@691 N_OUT9_Mn9@691_d N_OUT8_Mn9@691_g N_VSS_Mn9@691_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@690 N_OUT9_Mn9@690_d N_OUT8_Mn9@690_g N_VSS_Mn9@690_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@691 N_OUT9_Mp9@691_d N_OUT8_Mp9@691_g N_VDD_Mp9@691_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@690 N_OUT9_Mp9@690_d N_OUT8_Mp9@690_g N_VDD_Mp9@690_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@689 N_OUT9_Mn9@689_d N_OUT8_Mn9@689_g N_VSS_Mn9@689_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@688 N_OUT9_Mn9@688_d N_OUT8_Mn9@688_g N_VSS_Mn9@688_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@689 N_OUT9_Mp9@689_d N_OUT8_Mp9@689_g N_VDD_Mp9@689_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@688 N_OUT9_Mp9@688_d N_OUT8_Mp9@688_g N_VDD_Mp9@688_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@687 N_OUT9_Mn9@687_d N_OUT8_Mn9@687_g N_VSS_Mn9@687_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@686 N_OUT9_Mn9@686_d N_OUT8_Mn9@686_g N_VSS_Mn9@686_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@687 N_OUT9_Mp9@687_d N_OUT8_Mp9@687_g N_VDD_Mp9@687_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@686 N_OUT9_Mp9@686_d N_OUT8_Mp9@686_g N_VDD_Mp9@686_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@685 N_OUT9_Mn9@685_d N_OUT8_Mn9@685_g N_VSS_Mn9@685_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@684 N_OUT9_Mn9@684_d N_OUT8_Mn9@684_g N_VSS_Mn9@684_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@685 N_OUT9_Mp9@685_d N_OUT8_Mp9@685_g N_VDD_Mp9@685_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@684 N_OUT9_Mp9@684_d N_OUT8_Mp9@684_g N_VDD_Mp9@684_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@683 N_OUT9_Mn9@683_d N_OUT8_Mn9@683_g N_VSS_Mn9@683_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@682 N_OUT9_Mn9@682_d N_OUT8_Mn9@682_g N_VSS_Mn9@682_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@683 N_OUT9_Mp9@683_d N_OUT8_Mp9@683_g N_VDD_Mp9@683_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@682 N_OUT9_Mp9@682_d N_OUT8_Mp9@682_g N_VDD_Mp9@682_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@681 N_OUT9_Mn9@681_d N_OUT8_Mn9@681_g N_VSS_Mn9@681_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@680 N_OUT9_Mn9@680_d N_OUT8_Mn9@680_g N_VSS_Mn9@680_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@681 N_OUT9_Mp9@681_d N_OUT8_Mp9@681_g N_VDD_Mp9@681_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@680 N_OUT9_Mp9@680_d N_OUT8_Mp9@680_g N_VDD_Mp9@680_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@679 N_OUT9_Mn9@679_d N_OUT8_Mn9@679_g N_VSS_Mn9@679_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@678 N_OUT9_Mn9@678_d N_OUT8_Mn9@678_g N_VSS_Mn9@678_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@679 N_OUT9_Mp9@679_d N_OUT8_Mp9@679_g N_VDD_Mp9@679_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@678 N_OUT9_Mp9@678_d N_OUT8_Mp9@678_g N_VDD_Mp9@678_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@677 N_OUT9_Mn9@677_d N_OUT8_Mn9@677_g N_VSS_Mn9@677_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@676 N_OUT9_Mn9@676_d N_OUT8_Mn9@676_g N_VSS_Mn9@676_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@677 N_OUT9_Mp9@677_d N_OUT8_Mp9@677_g N_VDD_Mp9@677_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@676 N_OUT9_Mp9@676_d N_OUT8_Mp9@676_g N_VDD_Mp9@676_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@675 N_OUT9_Mn9@675_d N_OUT8_Mn9@675_g N_VSS_Mn9@675_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@674 N_OUT9_Mn9@674_d N_OUT8_Mn9@674_g N_VSS_Mn9@674_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@675 N_OUT9_Mp9@675_d N_OUT8_Mp9@675_g N_VDD_Mp9@675_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@674 N_OUT9_Mp9@674_d N_OUT8_Mp9@674_g N_VDD_Mp9@674_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@673 N_OUT9_Mn9@673_d N_OUT8_Mn9@673_g N_VSS_Mn9@673_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@672 N_OUT9_Mn9@672_d N_OUT8_Mn9@672_g N_VSS_Mn9@672_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@673 N_OUT9_Mp9@673_d N_OUT8_Mp9@673_g N_VDD_Mp9@673_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@672 N_OUT9_Mp9@672_d N_OUT8_Mp9@672_g N_VDD_Mp9@672_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@671 N_OUT9_Mn9@671_d N_OUT8_Mn9@671_g N_VSS_Mn9@671_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@670 N_OUT9_Mn9@670_d N_OUT8_Mn9@670_g N_VSS_Mn9@670_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@671 N_OUT9_Mp9@671_d N_OUT8_Mp9@671_g N_VDD_Mp9@671_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@670 N_OUT9_Mp9@670_d N_OUT8_Mp9@670_g N_VDD_Mp9@670_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@669 N_OUT9_Mn9@669_d N_OUT8_Mn9@669_g N_VSS_Mn9@669_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@668 N_OUT9_Mn9@668_d N_OUT8_Mn9@668_g N_VSS_Mn9@668_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@669 N_OUT9_Mp9@669_d N_OUT8_Mp9@669_g N_VDD_Mp9@669_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@668 N_OUT9_Mp9@668_d N_OUT8_Mp9@668_g N_VDD_Mp9@668_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@667 N_OUT9_Mn9@667_d N_OUT8_Mn9@667_g N_VSS_Mn9@667_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@666 N_OUT9_Mn9@666_d N_OUT8_Mn9@666_g N_VSS_Mn9@666_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@667 N_OUT9_Mp9@667_d N_OUT8_Mp9@667_g N_VDD_Mp9@667_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@666 N_OUT9_Mp9@666_d N_OUT8_Mp9@666_g N_VDD_Mp9@666_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@665 N_OUT9_Mn9@665_d N_OUT8_Mn9@665_g N_VSS_Mn9@665_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@664 N_OUT9_Mn9@664_d N_OUT8_Mn9@664_g N_VSS_Mn9@664_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@665 N_OUT9_Mp9@665_d N_OUT8_Mp9@665_g N_VDD_Mp9@665_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@664 N_OUT9_Mp9@664_d N_OUT8_Mp9@664_g N_VDD_Mp9@664_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@663 N_OUT9_Mn9@663_d N_OUT8_Mn9@663_g N_VSS_Mn9@663_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@662 N_OUT9_Mn9@662_d N_OUT8_Mn9@662_g N_VSS_Mn9@662_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@663 N_OUT9_Mp9@663_d N_OUT8_Mp9@663_g N_VDD_Mp9@663_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@662 N_OUT9_Mp9@662_d N_OUT8_Mp9@662_g N_VDD_Mp9@662_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@661 N_OUT9_Mn9@661_d N_OUT8_Mn9@661_g N_VSS_Mn9@661_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@660 N_OUT9_Mn9@660_d N_OUT8_Mn9@660_g N_VSS_Mn9@660_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@661 N_OUT9_Mp9@661_d N_OUT8_Mp9@661_g N_VDD_Mp9@661_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@660 N_OUT9_Mp9@660_d N_OUT8_Mp9@660_g N_VDD_Mp9@660_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@659 N_OUT9_Mn9@659_d N_OUT8_Mn9@659_g N_VSS_Mn9@659_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@658 N_OUT9_Mn9@658_d N_OUT8_Mn9@658_g N_VSS_Mn9@658_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@659 N_OUT9_Mp9@659_d N_OUT8_Mp9@659_g N_VDD_Mp9@659_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@658 N_OUT9_Mp9@658_d N_OUT8_Mp9@658_g N_VDD_Mp9@658_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@657 N_OUT9_Mn9@657_d N_OUT8_Mn9@657_g N_VSS_Mn9@657_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@656 N_OUT9_Mn9@656_d N_OUT8_Mn9@656_g N_VSS_Mn9@656_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@657 N_OUT9_Mp9@657_d N_OUT8_Mp9@657_g N_VDD_Mp9@657_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@656 N_OUT9_Mp9@656_d N_OUT8_Mp9@656_g N_VDD_Mp9@656_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@655 N_OUT9_Mn9@655_d N_OUT8_Mn9@655_g N_VSS_Mn9@655_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@654 N_OUT9_Mn9@654_d N_OUT8_Mn9@654_g N_VSS_Mn9@654_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@655 N_OUT9_Mp9@655_d N_OUT8_Mp9@655_g N_VDD_Mp9@655_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@654 N_OUT9_Mp9@654_d N_OUT8_Mp9@654_g N_VDD_Mp9@654_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@653 N_OUT9_Mn9@653_d N_OUT8_Mn9@653_g N_VSS_Mn9@653_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@652 N_OUT9_Mn9@652_d N_OUT8_Mn9@652_g N_VSS_Mn9@652_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@653 N_OUT9_Mp9@653_d N_OUT8_Mp9@653_g N_VDD_Mp9@653_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@652 N_OUT9_Mp9@652_d N_OUT8_Mp9@652_g N_VDD_Mp9@652_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@651 N_OUT9_Mn9@651_d N_OUT8_Mn9@651_g N_VSS_Mn9@651_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@650 N_OUT9_Mn9@650_d N_OUT8_Mn9@650_g N_VSS_Mn9@650_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@651 N_OUT9_Mp9@651_d N_OUT8_Mp9@651_g N_VDD_Mp9@651_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@650 N_OUT9_Mp9@650_d N_OUT8_Mp9@650_g N_VDD_Mp9@650_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@649 N_OUT9_Mn9@649_d N_OUT8_Mn9@649_g N_VSS_Mn9@649_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@648 N_OUT9_Mn9@648_d N_OUT8_Mn9@648_g N_VSS_Mn9@648_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@649 N_OUT9_Mp9@649_d N_OUT8_Mp9@649_g N_VDD_Mp9@649_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@648 N_OUT9_Mp9@648_d N_OUT8_Mp9@648_g N_VDD_Mp9@648_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@647 N_OUT9_Mn9@647_d N_OUT8_Mn9@647_g N_VSS_Mn9@647_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@646 N_OUT9_Mn9@646_d N_OUT8_Mn9@646_g N_VSS_Mn9@646_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@647 N_OUT9_Mp9@647_d N_OUT8_Mp9@647_g N_VDD_Mp9@647_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@646 N_OUT9_Mp9@646_d N_OUT8_Mp9@646_g N_VDD_Mp9@646_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@645 N_OUT9_Mn9@645_d N_OUT8_Mn9@645_g N_VSS_Mn9@645_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@644 N_OUT9_Mn9@644_d N_OUT8_Mn9@644_g N_VSS_Mn9@644_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@645 N_OUT9_Mp9@645_d N_OUT8_Mp9@645_g N_VDD_Mp9@645_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@644 N_OUT9_Mp9@644_d N_OUT8_Mp9@644_g N_VDD_Mp9@644_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@643 N_OUT9_Mn9@643_d N_OUT8_Mn9@643_g N_VSS_Mn9@643_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@642 N_OUT9_Mn9@642_d N_OUT8_Mn9@642_g N_VSS_Mn9@642_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@643 N_OUT9_Mp9@643_d N_OUT8_Mp9@643_g N_VDD_Mp9@643_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@642 N_OUT9_Mp9@642_d N_OUT8_Mp9@642_g N_VDD_Mp9@642_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@641 N_OUT9_Mn9@641_d N_OUT8_Mn9@641_g N_VSS_Mn9@641_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@640 N_OUT9_Mn9@640_d N_OUT8_Mn9@640_g N_VSS_Mn9@640_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@641 N_OUT9_Mp9@641_d N_OUT8_Mp9@641_g N_VDD_Mp9@641_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@640 N_OUT9_Mp9@640_d N_OUT8_Mp9@640_g N_VDD_Mp9@640_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@639 N_OUT9_Mn9@639_d N_OUT8_Mn9@639_g N_VSS_Mn9@639_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@638 N_OUT9_Mn9@638_d N_OUT8_Mn9@638_g N_VSS_Mn9@638_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@639 N_OUT9_Mp9@639_d N_OUT8_Mp9@639_g N_VDD_Mp9@639_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@638 N_OUT9_Mp9@638_d N_OUT8_Mp9@638_g N_VDD_Mp9@638_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@637 N_OUT9_Mn9@637_d N_OUT8_Mn9@637_g N_VSS_Mn9@637_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@636 N_OUT9_Mn9@636_d N_OUT8_Mn9@636_g N_VSS_Mn9@636_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@637 N_OUT9_Mp9@637_d N_OUT8_Mp9@637_g N_VDD_Mp9@637_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@636 N_OUT9_Mp9@636_d N_OUT8_Mp9@636_g N_VDD_Mp9@636_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@635 N_OUT9_Mn9@635_d N_OUT8_Mn9@635_g N_VSS_Mn9@635_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@634 N_OUT9_Mn9@634_d N_OUT8_Mn9@634_g N_VSS_Mn9@634_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@635 N_OUT9_Mp9@635_d N_OUT8_Mp9@635_g N_VDD_Mp9@635_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@634 N_OUT9_Mp9@634_d N_OUT8_Mp9@634_g N_VDD_Mp9@634_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@633 N_OUT9_Mn9@633_d N_OUT8_Mn9@633_g N_VSS_Mn9@633_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@632 N_OUT9_Mn9@632_d N_OUT8_Mn9@632_g N_VSS_Mn9@632_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@633 N_OUT9_Mp9@633_d N_OUT8_Mp9@633_g N_VDD_Mp9@633_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@632 N_OUT9_Mp9@632_d N_OUT8_Mp9@632_g N_VDD_Mp9@632_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@631 N_OUT9_Mn9@631_d N_OUT8_Mn9@631_g N_VSS_Mn9@631_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@630 N_OUT9_Mn9@630_d N_OUT8_Mn9@630_g N_VSS_Mn9@630_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@631 N_OUT9_Mp9@631_d N_OUT8_Mp9@631_g N_VDD_Mp9@631_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@630 N_OUT9_Mp9@630_d N_OUT8_Mp9@630_g N_VDD_Mp9@630_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@629 N_OUT9_Mn9@629_d N_OUT8_Mn9@629_g N_VSS_Mn9@629_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@628 N_OUT9_Mn9@628_d N_OUT8_Mn9@628_g N_VSS_Mn9@628_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@629 N_OUT9_Mp9@629_d N_OUT8_Mp9@629_g N_VDD_Mp9@629_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@628 N_OUT9_Mp9@628_d N_OUT8_Mp9@628_g N_VDD_Mp9@628_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@627 N_OUT9_Mn9@627_d N_OUT8_Mn9@627_g N_VSS_Mn9@627_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@626 N_OUT9_Mn9@626_d N_OUT8_Mn9@626_g N_VSS_Mn9@626_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@627 N_OUT9_Mp9@627_d N_OUT8_Mp9@627_g N_VDD_Mp9@627_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@626 N_OUT9_Mp9@626_d N_OUT8_Mp9@626_g N_VDD_Mp9@626_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@625 N_OUT9_Mn9@625_d N_OUT8_Mn9@625_g N_VSS_Mn9@625_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@624 N_OUT9_Mn9@624_d N_OUT8_Mn9@624_g N_VSS_Mn9@624_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@625 N_OUT9_Mp9@625_d N_OUT8_Mp9@625_g N_VDD_Mp9@625_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@624 N_OUT9_Mp9@624_d N_OUT8_Mp9@624_g N_VDD_Mp9@624_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@623 N_OUT9_Mn9@623_d N_OUT8_Mn9@623_g N_VSS_Mn9@623_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@622 N_OUT9_Mn9@622_d N_OUT8_Mn9@622_g N_VSS_Mn9@622_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@623 N_OUT9_Mp9@623_d N_OUT8_Mp9@623_g N_VDD_Mp9@623_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@622 N_OUT9_Mp9@622_d N_OUT8_Mp9@622_g N_VDD_Mp9@622_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@621 N_OUT9_Mn9@621_d N_OUT8_Mn9@621_g N_VSS_Mn9@621_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@620 N_OUT9_Mn9@620_d N_OUT8_Mn9@620_g N_VSS_Mn9@620_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@621 N_OUT9_Mp9@621_d N_OUT8_Mp9@621_g N_VDD_Mp9@621_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@620 N_OUT9_Mp9@620_d N_OUT8_Mp9@620_g N_VDD_Mp9@620_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@619 N_OUT9_Mn9@619_d N_OUT8_Mn9@619_g N_VSS_Mn9@619_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@618 N_OUT9_Mn9@618_d N_OUT8_Mn9@618_g N_VSS_Mn9@618_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@619 N_OUT9_Mp9@619_d N_OUT8_Mp9@619_g N_VDD_Mp9@619_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@618 N_OUT9_Mp9@618_d N_OUT8_Mp9@618_g N_VDD_Mp9@618_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@617 N_OUT9_Mn9@617_d N_OUT8_Mn9@617_g N_VSS_Mn9@617_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@616 N_OUT9_Mn9@616_d N_OUT8_Mn9@616_g N_VSS_Mn9@616_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@617 N_OUT9_Mp9@617_d N_OUT8_Mp9@617_g N_VDD_Mp9@617_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@616 N_OUT9_Mp9@616_d N_OUT8_Mp9@616_g N_VDD_Mp9@616_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@615 N_OUT9_Mn9@615_d N_OUT8_Mn9@615_g N_VSS_Mn9@615_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@614 N_OUT9_Mn9@614_d N_OUT8_Mn9@614_g N_VSS_Mn9@614_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@615 N_OUT9_Mp9@615_d N_OUT8_Mp9@615_g N_VDD_Mp9@615_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@614 N_OUT9_Mp9@614_d N_OUT8_Mp9@614_g N_VDD_Mp9@614_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@613 N_OUT9_Mn9@613_d N_OUT8_Mn9@613_g N_VSS_Mn9@613_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@612 N_OUT9_Mn9@612_d N_OUT8_Mn9@612_g N_VSS_Mn9@612_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@613 N_OUT9_Mp9@613_d N_OUT8_Mp9@613_g N_VDD_Mp9@613_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@612 N_OUT9_Mp9@612_d N_OUT8_Mp9@612_g N_VDD_Mp9@612_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@611 N_OUT9_Mn9@611_d N_OUT8_Mn9@611_g N_VSS_Mn9@611_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@610 N_OUT9_Mn9@610_d N_OUT8_Mn9@610_g N_VSS_Mn9@610_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@611 N_OUT9_Mp9@611_d N_OUT8_Mp9@611_g N_VDD_Mp9@611_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@610 N_OUT9_Mp9@610_d N_OUT8_Mp9@610_g N_VDD_Mp9@610_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@609 N_OUT9_Mn9@609_d N_OUT8_Mn9@609_g N_VSS_Mn9@609_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@608 N_OUT9_Mn9@608_d N_OUT8_Mn9@608_g N_VSS_Mn9@608_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@609 N_OUT9_Mp9@609_d N_OUT8_Mp9@609_g N_VDD_Mp9@609_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@608 N_OUT9_Mp9@608_d N_OUT8_Mp9@608_g N_VDD_Mp9@608_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@607 N_OUT9_Mn9@607_d N_OUT8_Mn9@607_g N_VSS_Mn9@607_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@606 N_OUT9_Mn9@606_d N_OUT8_Mn9@606_g N_VSS_Mn9@606_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@607 N_OUT9_Mp9@607_d N_OUT8_Mp9@607_g N_VDD_Mp9@607_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@606 N_OUT9_Mp9@606_d N_OUT8_Mp9@606_g N_VDD_Mp9@606_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@605 N_OUT9_Mn9@605_d N_OUT8_Mn9@605_g N_VSS_Mn9@605_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@604 N_OUT9_Mn9@604_d N_OUT8_Mn9@604_g N_VSS_Mn9@604_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@605 N_OUT9_Mp9@605_d N_OUT8_Mp9@605_g N_VDD_Mp9@605_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@604 N_OUT9_Mp9@604_d N_OUT8_Mp9@604_g N_VDD_Mp9@604_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@603 N_OUT9_Mn9@603_d N_OUT8_Mn9@603_g N_VSS_Mn9@603_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@602 N_OUT9_Mn9@602_d N_OUT8_Mn9@602_g N_VSS_Mn9@602_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@603 N_OUT9_Mp9@603_d N_OUT8_Mp9@603_g N_VDD_Mp9@603_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@602 N_OUT9_Mp9@602_d N_OUT8_Mp9@602_g N_VDD_Mp9@602_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@601 N_OUT9_Mn9@601_d N_OUT8_Mn9@601_g N_VSS_Mn9@601_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@600 N_OUT9_Mn9@600_d N_OUT8_Mn9@600_g N_VSS_Mn9@600_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@601 N_OUT9_Mp9@601_d N_OUT8_Mp9@601_g N_VDD_Mp9@601_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@600 N_OUT9_Mp9@600_d N_OUT8_Mp9@600_g N_VDD_Mp9@600_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@599 N_OUT9_Mn9@599_d N_OUT8_Mn9@599_g N_VSS_Mn9@599_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@598 N_OUT9_Mn9@598_d N_OUT8_Mn9@598_g N_VSS_Mn9@598_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@599 N_OUT9_Mp9@599_d N_OUT8_Mp9@599_g N_VDD_Mp9@599_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@598 N_OUT9_Mp9@598_d N_OUT8_Mp9@598_g N_VDD_Mp9@598_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@597 N_OUT9_Mn9@597_d N_OUT8_Mn9@597_g N_VSS_Mn9@597_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@596 N_OUT9_Mn9@596_d N_OUT8_Mn9@596_g N_VSS_Mn9@596_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@597 N_OUT9_Mp9@597_d N_OUT8_Mp9@597_g N_VDD_Mp9@597_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@596 N_OUT9_Mp9@596_d N_OUT8_Mp9@596_g N_VDD_Mp9@596_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@595 N_OUT9_Mn9@595_d N_OUT8_Mn9@595_g N_VSS_Mn9@595_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@594 N_OUT9_Mn9@594_d N_OUT8_Mn9@594_g N_VSS_Mn9@594_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@595 N_OUT9_Mp9@595_d N_OUT8_Mp9@595_g N_VDD_Mp9@595_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@594 N_OUT9_Mp9@594_d N_OUT8_Mp9@594_g N_VDD_Mp9@594_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@593 N_OUT9_Mn9@593_d N_OUT8_Mn9@593_g N_VSS_Mn9@593_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@592 N_OUT9_Mn9@592_d N_OUT8_Mn9@592_g N_VSS_Mn9@592_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@593 N_OUT9_Mp9@593_d N_OUT8_Mp9@593_g N_VDD_Mp9@593_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@592 N_OUT9_Mp9@592_d N_OUT8_Mp9@592_g N_VDD_Mp9@592_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@591 N_OUT9_Mn9@591_d N_OUT8_Mn9@591_g N_VSS_Mn9@591_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@590 N_OUT9_Mn9@590_d N_OUT8_Mn9@590_g N_VSS_Mn9@590_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@591 N_OUT9_Mp9@591_d N_OUT8_Mp9@591_g N_VDD_Mp9@591_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@590 N_OUT9_Mp9@590_d N_OUT8_Mp9@590_g N_VDD_Mp9@590_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@589 N_OUT9_Mn9@589_d N_OUT8_Mn9@589_g N_VSS_Mn9@589_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@588 N_OUT9_Mn9@588_d N_OUT8_Mn9@588_g N_VSS_Mn9@588_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@589 N_OUT9_Mp9@589_d N_OUT8_Mp9@589_g N_VDD_Mp9@589_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@588 N_OUT9_Mp9@588_d N_OUT8_Mp9@588_g N_VDD_Mp9@588_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@587 N_OUT9_Mn9@587_d N_OUT8_Mn9@587_g N_VSS_Mn9@587_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@586 N_OUT9_Mn9@586_d N_OUT8_Mn9@586_g N_VSS_Mn9@586_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@587 N_OUT9_Mp9@587_d N_OUT8_Mp9@587_g N_VDD_Mp9@587_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@586 N_OUT9_Mp9@586_d N_OUT8_Mp9@586_g N_VDD_Mp9@586_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@585 N_OUT9_Mn9@585_d N_OUT8_Mn9@585_g N_VSS_Mn9@585_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@584 N_OUT9_Mn9@584_d N_OUT8_Mn9@584_g N_VSS_Mn9@584_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@585 N_OUT9_Mp9@585_d N_OUT8_Mp9@585_g N_VDD_Mp9@585_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@584 N_OUT9_Mp9@584_d N_OUT8_Mp9@584_g N_VDD_Mp9@584_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@583 N_OUT9_Mn9@583_d N_OUT8_Mn9@583_g N_VSS_Mn9@583_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@582 N_OUT9_Mn9@582_d N_OUT8_Mn9@582_g N_VSS_Mn9@582_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@583 N_OUT9_Mp9@583_d N_OUT8_Mp9@583_g N_VDD_Mp9@583_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@582 N_OUT9_Mp9@582_d N_OUT8_Mp9@582_g N_VDD_Mp9@582_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@581 N_OUT9_Mn9@581_d N_OUT8_Mn9@581_g N_VSS_Mn9@581_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@580 N_OUT9_Mn9@580_d N_OUT8_Mn9@580_g N_VSS_Mn9@580_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@581 N_OUT9_Mp9@581_d N_OUT8_Mp9@581_g N_VDD_Mp9@581_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@580 N_OUT9_Mp9@580_d N_OUT8_Mp9@580_g N_VDD_Mp9@580_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@579 N_OUT9_Mn9@579_d N_OUT8_Mn9@579_g N_VSS_Mn9@579_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@578 N_OUT9_Mn9@578_d N_OUT8_Mn9@578_g N_VSS_Mn9@578_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@579 N_OUT9_Mp9@579_d N_OUT8_Mp9@579_g N_VDD_Mp9@579_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@578 N_OUT9_Mp9@578_d N_OUT8_Mp9@578_g N_VDD_Mp9@578_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@577 N_OUT9_Mn9@577_d N_OUT8_Mn9@577_g N_VSS_Mn9@577_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@576 N_OUT9_Mn9@576_d N_OUT8_Mn9@576_g N_VSS_Mn9@576_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@577 N_OUT9_Mp9@577_d N_OUT8_Mp9@577_g N_VDD_Mp9@577_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@576 N_OUT9_Mp9@576_d N_OUT8_Mp9@576_g N_VDD_Mp9@576_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@575 N_OUT9_Mn9@575_d N_OUT8_Mn9@575_g N_VSS_Mn9@575_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@574 N_OUT9_Mn9@574_d N_OUT8_Mn9@574_g N_VSS_Mn9@574_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@575 N_OUT9_Mp9@575_d N_OUT8_Mp9@575_g N_VDD_Mp9@575_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@574 N_OUT9_Mp9@574_d N_OUT8_Mp9@574_g N_VDD_Mp9@574_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@573 N_OUT9_Mn9@573_d N_OUT8_Mn9@573_g N_VSS_Mn9@573_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@572 N_OUT9_Mn9@572_d N_OUT8_Mn9@572_g N_VSS_Mn9@572_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@573 N_OUT9_Mp9@573_d N_OUT8_Mp9@573_g N_VDD_Mp9@573_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@572 N_OUT9_Mp9@572_d N_OUT8_Mp9@572_g N_VDD_Mp9@572_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@571 N_OUT9_Mn9@571_d N_OUT8_Mn9@571_g N_VSS_Mn9@571_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@570 N_OUT9_Mn9@570_d N_OUT8_Mn9@570_g N_VSS_Mn9@570_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@571 N_OUT9_Mp9@571_d N_OUT8_Mp9@571_g N_VDD_Mp9@571_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@570 N_OUT9_Mp9@570_d N_OUT8_Mp9@570_g N_VDD_Mp9@570_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@569 N_OUT9_Mn9@569_d N_OUT8_Mn9@569_g N_VSS_Mn9@569_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@568 N_OUT9_Mn9@568_d N_OUT8_Mn9@568_g N_VSS_Mn9@568_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@569 N_OUT9_Mp9@569_d N_OUT8_Mp9@569_g N_VDD_Mp9@569_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@568 N_OUT9_Mp9@568_d N_OUT8_Mp9@568_g N_VDD_Mp9@568_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@567 N_OUT9_Mn9@567_d N_OUT8_Mn9@567_g N_VSS_Mn9@567_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@566 N_OUT9_Mn9@566_d N_OUT8_Mn9@566_g N_VSS_Mn9@566_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@567 N_OUT9_Mp9@567_d N_OUT8_Mp9@567_g N_VDD_Mp9@567_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@566 N_OUT9_Mp9@566_d N_OUT8_Mp9@566_g N_VDD_Mp9@566_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@565 N_OUT9_Mn9@565_d N_OUT8_Mn9@565_g N_VSS_Mn9@565_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@564 N_OUT9_Mn9@564_d N_OUT8_Mn9@564_g N_VSS_Mn9@564_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@565 N_OUT9_Mp9@565_d N_OUT8_Mp9@565_g N_VDD_Mp9@565_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@564 N_OUT9_Mp9@564_d N_OUT8_Mp9@564_g N_VDD_Mp9@564_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@563 N_OUT9_Mn9@563_d N_OUT8_Mn9@563_g N_VSS_Mn9@563_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@562 N_OUT9_Mn9@562_d N_OUT8_Mn9@562_g N_VSS_Mn9@562_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@563 N_OUT9_Mp9@563_d N_OUT8_Mp9@563_g N_VDD_Mp9@563_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@562 N_OUT9_Mp9@562_d N_OUT8_Mp9@562_g N_VDD_Mp9@562_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@561 N_OUT9_Mn9@561_d N_OUT8_Mn9@561_g N_VSS_Mn9@561_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@560 N_OUT9_Mn9@560_d N_OUT8_Mn9@560_g N_VSS_Mn9@560_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@561 N_OUT9_Mp9@561_d N_OUT8_Mp9@561_g N_VDD_Mp9@561_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@560 N_OUT9_Mp9@560_d N_OUT8_Mp9@560_g N_VDD_Mp9@560_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@559 N_OUT9_Mn9@559_d N_OUT8_Mn9@559_g N_VSS_Mn9@559_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@558 N_OUT9_Mn9@558_d N_OUT8_Mn9@558_g N_VSS_Mn9@558_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@559 N_OUT9_Mp9@559_d N_OUT8_Mp9@559_g N_VDD_Mp9@559_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@558 N_OUT9_Mp9@558_d N_OUT8_Mp9@558_g N_VDD_Mp9@558_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@557 N_OUT9_Mn9@557_d N_OUT8_Mn9@557_g N_VSS_Mn9@557_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@556 N_OUT9_Mn9@556_d N_OUT8_Mn9@556_g N_VSS_Mn9@556_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@557 N_OUT9_Mp9@557_d N_OUT8_Mp9@557_g N_VDD_Mp9@557_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@556 N_OUT9_Mp9@556_d N_OUT8_Mp9@556_g N_VDD_Mp9@556_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@555 N_OUT9_Mn9@555_d N_OUT8_Mn9@555_g N_VSS_Mn9@555_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@554 N_OUT9_Mn9@554_d N_OUT8_Mn9@554_g N_VSS_Mn9@554_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@555 N_OUT9_Mp9@555_d N_OUT8_Mp9@555_g N_VDD_Mp9@555_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@554 N_OUT9_Mp9@554_d N_OUT8_Mp9@554_g N_VDD_Mp9@554_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@553 N_OUT9_Mn9@553_d N_OUT8_Mn9@553_g N_VSS_Mn9@553_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@552 N_OUT9_Mn9@552_d N_OUT8_Mn9@552_g N_VSS_Mn9@552_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@553 N_OUT9_Mp9@553_d N_OUT8_Mp9@553_g N_VDD_Mp9@553_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@552 N_OUT9_Mp9@552_d N_OUT8_Mp9@552_g N_VDD_Mp9@552_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@551 N_OUT9_Mn9@551_d N_OUT8_Mn9@551_g N_VSS_Mn9@551_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@550 N_OUT9_Mn9@550_d N_OUT8_Mn9@550_g N_VSS_Mn9@550_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@551 N_OUT9_Mp9@551_d N_OUT8_Mp9@551_g N_VDD_Mp9@551_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@550 N_OUT9_Mp9@550_d N_OUT8_Mp9@550_g N_VDD_Mp9@550_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@549 N_OUT9_Mn9@549_d N_OUT8_Mn9@549_g N_VSS_Mn9@549_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@548 N_OUT9_Mn9@548_d N_OUT8_Mn9@548_g N_VSS_Mn9@548_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@549 N_OUT9_Mp9@549_d N_OUT8_Mp9@549_g N_VDD_Mp9@549_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@548 N_OUT9_Mp9@548_d N_OUT8_Mp9@548_g N_VDD_Mp9@548_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@547 N_OUT9_Mn9@547_d N_OUT8_Mn9@547_g N_VSS_Mn9@547_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@546 N_OUT9_Mn9@546_d N_OUT8_Mn9@546_g N_VSS_Mn9@546_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@547 N_OUT9_Mp9@547_d N_OUT8_Mp9@547_g N_VDD_Mp9@547_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@546 N_OUT9_Mp9@546_d N_OUT8_Mp9@546_g N_VDD_Mp9@546_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@545 N_OUT9_Mn9@545_d N_OUT8_Mn9@545_g N_VSS_Mn9@545_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@544 N_OUT9_Mn9@544_d N_OUT8_Mn9@544_g N_VSS_Mn9@544_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@545 N_OUT9_Mp9@545_d N_OUT8_Mp9@545_g N_VDD_Mp9@545_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@544 N_OUT9_Mp9@544_d N_OUT8_Mp9@544_g N_VDD_Mp9@544_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@543 N_OUT9_Mn9@543_d N_OUT8_Mn9@543_g N_VSS_Mn9@543_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@542 N_OUT9_Mn9@542_d N_OUT8_Mn9@542_g N_VSS_Mn9@542_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@543 N_OUT9_Mp9@543_d N_OUT8_Mp9@543_g N_VDD_Mp9@543_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@542 N_OUT9_Mp9@542_d N_OUT8_Mp9@542_g N_VDD_Mp9@542_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@541 N_OUT9_Mn9@541_d N_OUT8_Mn9@541_g N_VSS_Mn9@541_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@540 N_OUT9_Mn9@540_d N_OUT8_Mn9@540_g N_VSS_Mn9@540_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@541 N_OUT9_Mp9@541_d N_OUT8_Mp9@541_g N_VDD_Mp9@541_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@540 N_OUT9_Mp9@540_d N_OUT8_Mp9@540_g N_VDD_Mp9@540_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@539 N_OUT9_Mn9@539_d N_OUT8_Mn9@539_g N_VSS_Mn9@539_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@538 N_OUT9_Mn9@538_d N_OUT8_Mn9@538_g N_VSS_Mn9@538_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@539 N_OUT9_Mp9@539_d N_OUT8_Mp9@539_g N_VDD_Mp9@539_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@538 N_OUT9_Mp9@538_d N_OUT8_Mp9@538_g N_VDD_Mp9@538_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@537 N_OUT9_Mn9@537_d N_OUT8_Mn9@537_g N_VSS_Mn9@537_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@536 N_OUT9_Mn9@536_d N_OUT8_Mn9@536_g N_VSS_Mn9@536_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@537 N_OUT9_Mp9@537_d N_OUT8_Mp9@537_g N_VDD_Mp9@537_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@536 N_OUT9_Mp9@536_d N_OUT8_Mp9@536_g N_VDD_Mp9@536_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@535 N_OUT9_Mn9@535_d N_OUT8_Mn9@535_g N_VSS_Mn9@535_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@534 N_OUT9_Mn9@534_d N_OUT8_Mn9@534_g N_VSS_Mn9@534_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@535 N_OUT9_Mp9@535_d N_OUT8_Mp9@535_g N_VDD_Mp9@535_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@534 N_OUT9_Mp9@534_d N_OUT8_Mp9@534_g N_VDD_Mp9@534_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@533 N_OUT9_Mn9@533_d N_OUT8_Mn9@533_g N_VSS_Mn9@533_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@532 N_OUT9_Mn9@532_d N_OUT8_Mn9@532_g N_VSS_Mn9@532_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@533 N_OUT9_Mp9@533_d N_OUT8_Mp9@533_g N_VDD_Mp9@533_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@532 N_OUT9_Mp9@532_d N_OUT8_Mp9@532_g N_VDD_Mp9@532_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@531 N_OUT9_Mn9@531_d N_OUT8_Mn9@531_g N_VSS_Mn9@531_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@530 N_OUT9_Mn9@530_d N_OUT8_Mn9@530_g N_VSS_Mn9@530_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@531 N_OUT9_Mp9@531_d N_OUT8_Mp9@531_g N_VDD_Mp9@531_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@530 N_OUT9_Mp9@530_d N_OUT8_Mp9@530_g N_VDD_Mp9@530_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@529 N_OUT9_Mn9@529_d N_OUT8_Mn9@529_g N_VSS_Mn9@529_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@528 N_OUT9_Mn9@528_d N_OUT8_Mn9@528_g N_VSS_Mn9@528_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@529 N_OUT9_Mp9@529_d N_OUT8_Mp9@529_g N_VDD_Mp9@529_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@528 N_OUT9_Mp9@528_d N_OUT8_Mp9@528_g N_VDD_Mp9@528_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@527 N_OUT9_Mn9@527_d N_OUT8_Mn9@527_g N_VSS_Mn9@527_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@526 N_OUT9_Mn9@526_d N_OUT8_Mn9@526_g N_VSS_Mn9@526_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@527 N_OUT9_Mp9@527_d N_OUT8_Mp9@527_g N_VDD_Mp9@527_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@526 N_OUT9_Mp9@526_d N_OUT8_Mp9@526_g N_VDD_Mp9@526_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@525 N_OUT9_Mn9@525_d N_OUT8_Mn9@525_g N_VSS_Mn9@525_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@524 N_OUT9_Mn9@524_d N_OUT8_Mn9@524_g N_VSS_Mn9@524_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@525 N_OUT9_Mp9@525_d N_OUT8_Mp9@525_g N_VDD_Mp9@525_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@524 N_OUT9_Mp9@524_d N_OUT8_Mp9@524_g N_VDD_Mp9@524_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@523 N_OUT9_Mn9@523_d N_OUT8_Mn9@523_g N_VSS_Mn9@523_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@522 N_OUT9_Mn9@522_d N_OUT8_Mn9@522_g N_VSS_Mn9@522_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@523 N_OUT9_Mp9@523_d N_OUT8_Mp9@523_g N_VDD_Mp9@523_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@522 N_OUT9_Mp9@522_d N_OUT8_Mp9@522_g N_VDD_Mp9@522_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@521 N_OUT9_Mn9@521_d N_OUT8_Mn9@521_g N_VSS_Mn9@521_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@520 N_OUT9_Mn9@520_d N_OUT8_Mn9@520_g N_VSS_Mn9@520_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@521 N_OUT9_Mp9@521_d N_OUT8_Mp9@521_g N_VDD_Mp9@521_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@520 N_OUT9_Mp9@520_d N_OUT8_Mp9@520_g N_VDD_Mp9@520_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@519 N_OUT9_Mn9@519_d N_OUT8_Mn9@519_g N_VSS_Mn9@519_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@518 N_OUT9_Mn9@518_d N_OUT8_Mn9@518_g N_VSS_Mn9@518_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@519 N_OUT9_Mp9@519_d N_OUT8_Mp9@519_g N_VDD_Mp9@519_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@518 N_OUT9_Mp9@518_d N_OUT8_Mp9@518_g N_VDD_Mp9@518_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@517 N_OUT9_Mn9@517_d N_OUT8_Mn9@517_g N_VSS_Mn9@517_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@516 N_OUT9_Mn9@516_d N_OUT8_Mn9@516_g N_VSS_Mn9@516_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@517 N_OUT9_Mp9@517_d N_OUT8_Mp9@517_g N_VDD_Mp9@517_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@516 N_OUT9_Mp9@516_d N_OUT8_Mp9@516_g N_VDD_Mp9@516_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@515 N_OUT9_Mn9@515_d N_OUT8_Mn9@515_g N_VSS_Mn9@515_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@514 N_OUT9_Mn9@514_d N_OUT8_Mn9@514_g N_VSS_Mn9@514_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@515 N_OUT9_Mp9@515_d N_OUT8_Mp9@515_g N_VDD_Mp9@515_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@514 N_OUT9_Mp9@514_d N_OUT8_Mp9@514_g N_VDD_Mp9@514_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@513 N_OUT9_Mn9@513_d N_OUT8_Mn9@513_g N_VSS_Mn9@513_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@512 N_OUT9_Mn9@512_d N_OUT8_Mn9@512_g N_VSS_Mn9@512_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@513 N_OUT9_Mp9@513_d N_OUT8_Mp9@513_g N_VDD_Mp9@513_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@512 N_OUT9_Mp9@512_d N_OUT8_Mp9@512_g N_VDD_Mp9@512_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@511 N_OUT9_Mn9@511_d N_OUT8_Mn9@511_g N_VSS_Mn9@511_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@510 N_OUT9_Mn9@510_d N_OUT8_Mn9@510_g N_VSS_Mn9@510_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@511 N_OUT9_Mp9@511_d N_OUT8_Mp9@511_g N_VDD_Mp9@511_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@510 N_OUT9_Mp9@510_d N_OUT8_Mp9@510_g N_VDD_Mp9@510_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@509 N_OUT9_Mn9@509_d N_OUT8_Mn9@509_g N_VSS_Mn9@509_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@508 N_OUT9_Mn9@508_d N_OUT8_Mn9@508_g N_VSS_Mn9@508_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@509 N_OUT9_Mp9@509_d N_OUT8_Mp9@509_g N_VDD_Mp9@509_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@508 N_OUT9_Mp9@508_d N_OUT8_Mp9@508_g N_VDD_Mp9@508_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@507 N_OUT9_Mn9@507_d N_OUT8_Mn9@507_g N_VSS_Mn9@507_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@506 N_OUT9_Mn9@506_d N_OUT8_Mn9@506_g N_VSS_Mn9@506_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@507 N_OUT9_Mp9@507_d N_OUT8_Mp9@507_g N_VDD_Mp9@507_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@506 N_OUT9_Mp9@506_d N_OUT8_Mp9@506_g N_VDD_Mp9@506_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@505 N_OUT9_Mn9@505_d N_OUT8_Mn9@505_g N_VSS_Mn9@505_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@504 N_OUT9_Mn9@504_d N_OUT8_Mn9@504_g N_VSS_Mn9@504_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@505 N_OUT9_Mp9@505_d N_OUT8_Mp9@505_g N_VDD_Mp9@505_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@504 N_OUT9_Mp9@504_d N_OUT8_Mp9@504_g N_VDD_Mp9@504_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@503 N_OUT9_Mn9@503_d N_OUT8_Mn9@503_g N_VSS_Mn9@503_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@502 N_OUT9_Mn9@502_d N_OUT8_Mn9@502_g N_VSS_Mn9@502_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@503 N_OUT9_Mp9@503_d N_OUT8_Mp9@503_g N_VDD_Mp9@503_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@502 N_OUT9_Mp9@502_d N_OUT8_Mp9@502_g N_VDD_Mp9@502_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@501 N_OUT9_Mn9@501_d N_OUT8_Mn9@501_g N_VSS_Mn9@501_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@500 N_OUT9_Mn9@500_d N_OUT8_Mn9@500_g N_VSS_Mn9@500_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@501 N_OUT9_Mp9@501_d N_OUT8_Mp9@501_g N_VDD_Mp9@501_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@500 N_OUT9_Mp9@500_d N_OUT8_Mp9@500_g N_VDD_Mp9@500_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@499 N_OUT9_Mn9@499_d N_OUT8_Mn9@499_g N_VSS_Mn9@499_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@498 N_OUT9_Mn9@498_d N_OUT8_Mn9@498_g N_VSS_Mn9@498_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@499 N_OUT9_Mp9@499_d N_OUT8_Mp9@499_g N_VDD_Mp9@499_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@498 N_OUT9_Mp9@498_d N_OUT8_Mp9@498_g N_VDD_Mp9@498_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@497 N_OUT9_Mn9@497_d N_OUT8_Mn9@497_g N_VSS_Mn9@497_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@496 N_OUT9_Mn9@496_d N_OUT8_Mn9@496_g N_VSS_Mn9@496_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@497 N_OUT9_Mp9@497_d N_OUT8_Mp9@497_g N_VDD_Mp9@497_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@496 N_OUT9_Mp9@496_d N_OUT8_Mp9@496_g N_VDD_Mp9@496_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@495 N_OUT9_Mn9@495_d N_OUT8_Mn9@495_g N_VSS_Mn9@495_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@494 N_OUT9_Mn9@494_d N_OUT8_Mn9@494_g N_VSS_Mn9@494_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@495 N_OUT9_Mp9@495_d N_OUT8_Mp9@495_g N_VDD_Mp9@495_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@494 N_OUT9_Mp9@494_d N_OUT8_Mp9@494_g N_VDD_Mp9@494_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@493 N_OUT9_Mn9@493_d N_OUT8_Mn9@493_g N_VSS_Mn9@493_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@492 N_OUT9_Mn9@492_d N_OUT8_Mn9@492_g N_VSS_Mn9@492_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@493 N_OUT9_Mp9@493_d N_OUT8_Mp9@493_g N_VDD_Mp9@493_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@492 N_OUT9_Mp9@492_d N_OUT8_Mp9@492_g N_VDD_Mp9@492_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@491 N_OUT9_Mn9@491_d N_OUT8_Mn9@491_g N_VSS_Mn9@491_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@490 N_OUT9_Mn9@490_d N_OUT8_Mn9@490_g N_VSS_Mn9@490_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@491 N_OUT9_Mp9@491_d N_OUT8_Mp9@491_g N_VDD_Mp9@491_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@490 N_OUT9_Mp9@490_d N_OUT8_Mp9@490_g N_VDD_Mp9@490_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@489 N_OUT9_Mn9@489_d N_OUT8_Mn9@489_g N_VSS_Mn9@489_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@488 N_OUT9_Mn9@488_d N_OUT8_Mn9@488_g N_VSS_Mn9@488_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@489 N_OUT9_Mp9@489_d N_OUT8_Mp9@489_g N_VDD_Mp9@489_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@488 N_OUT9_Mp9@488_d N_OUT8_Mp9@488_g N_VDD_Mp9@488_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@487 N_OUT9_Mn9@487_d N_OUT8_Mn9@487_g N_VSS_Mn9@487_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@486 N_OUT9_Mn9@486_d N_OUT8_Mn9@486_g N_VSS_Mn9@486_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@487 N_OUT9_Mp9@487_d N_OUT8_Mp9@487_g N_VDD_Mp9@487_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@486 N_OUT9_Mp9@486_d N_OUT8_Mp9@486_g N_VDD_Mp9@486_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@485 N_OUT9_Mn9@485_d N_OUT8_Mn9@485_g N_VSS_Mn9@485_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@484 N_OUT9_Mn9@484_d N_OUT8_Mn9@484_g N_VSS_Mn9@484_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@485 N_OUT9_Mp9@485_d N_OUT8_Mp9@485_g N_VDD_Mp9@485_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@484 N_OUT9_Mp9@484_d N_OUT8_Mp9@484_g N_VDD_Mp9@484_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@483 N_OUT9_Mn9@483_d N_OUT8_Mn9@483_g N_VSS_Mn9@483_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@482 N_OUT9_Mn9@482_d N_OUT8_Mn9@482_g N_VSS_Mn9@482_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@483 N_OUT9_Mp9@483_d N_OUT8_Mp9@483_g N_VDD_Mp9@483_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@482 N_OUT9_Mp9@482_d N_OUT8_Mp9@482_g N_VDD_Mp9@482_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@481 N_OUT9_Mn9@481_d N_OUT8_Mn9@481_g N_VSS_Mn9@481_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@480 N_OUT9_Mn9@480_d N_OUT8_Mn9@480_g N_VSS_Mn9@480_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@481 N_OUT9_Mp9@481_d N_OUT8_Mp9@481_g N_VDD_Mp9@481_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@480 N_OUT9_Mp9@480_d N_OUT8_Mp9@480_g N_VDD_Mp9@480_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@479 N_OUT9_Mn9@479_d N_OUT8_Mn9@479_g N_VSS_Mn9@479_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@478 N_OUT9_Mn9@478_d N_OUT8_Mn9@478_g N_VSS_Mn9@478_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@479 N_OUT9_Mp9@479_d N_OUT8_Mp9@479_g N_VDD_Mp9@479_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@478 N_OUT9_Mp9@478_d N_OUT8_Mp9@478_g N_VDD_Mp9@478_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@477 N_OUT9_Mn9@477_d N_OUT8_Mn9@477_g N_VSS_Mn9@477_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@476 N_OUT9_Mn9@476_d N_OUT8_Mn9@476_g N_VSS_Mn9@476_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@477 N_OUT9_Mp9@477_d N_OUT8_Mp9@477_g N_VDD_Mp9@477_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@476 N_OUT9_Mp9@476_d N_OUT8_Mp9@476_g N_VDD_Mp9@476_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@475 N_OUT9_Mn9@475_d N_OUT8_Mn9@475_g N_VSS_Mn9@475_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@474 N_OUT9_Mn9@474_d N_OUT8_Mn9@474_g N_VSS_Mn9@474_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@475 N_OUT9_Mp9@475_d N_OUT8_Mp9@475_g N_VDD_Mp9@475_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@474 N_OUT9_Mp9@474_d N_OUT8_Mp9@474_g N_VDD_Mp9@474_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@473 N_OUT9_Mn9@473_d N_OUT8_Mn9@473_g N_VSS_Mn9@473_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@472 N_OUT9_Mn9@472_d N_OUT8_Mn9@472_g N_VSS_Mn9@472_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@473 N_OUT9_Mp9@473_d N_OUT8_Mp9@473_g N_VDD_Mp9@473_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@472 N_OUT9_Mp9@472_d N_OUT8_Mp9@472_g N_VDD_Mp9@472_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@471 N_OUT9_Mn9@471_d N_OUT8_Mn9@471_g N_VSS_Mn9@471_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@470 N_OUT9_Mn9@470_d N_OUT8_Mn9@470_g N_VSS_Mn9@470_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@471 N_OUT9_Mp9@471_d N_OUT8_Mp9@471_g N_VDD_Mp9@471_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@470 N_OUT9_Mp9@470_d N_OUT8_Mp9@470_g N_VDD_Mp9@470_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@469 N_OUT9_Mn9@469_d N_OUT8_Mn9@469_g N_VSS_Mn9@469_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@468 N_OUT9_Mn9@468_d N_OUT8_Mn9@468_g N_VSS_Mn9@468_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@469 N_OUT9_Mp9@469_d N_OUT8_Mp9@469_g N_VDD_Mp9@469_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@468 N_OUT9_Mp9@468_d N_OUT8_Mp9@468_g N_VDD_Mp9@468_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@467 N_OUT9_Mn9@467_d N_OUT8_Mn9@467_g N_VSS_Mn9@467_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@466 N_OUT9_Mn9@466_d N_OUT8_Mn9@466_g N_VSS_Mn9@466_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@467 N_OUT9_Mp9@467_d N_OUT8_Mp9@467_g N_VDD_Mp9@467_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@466 N_OUT9_Mp9@466_d N_OUT8_Mp9@466_g N_VDD_Mp9@466_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@465 N_OUT9_Mn9@465_d N_OUT8_Mn9@465_g N_VSS_Mn9@465_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@464 N_OUT9_Mn9@464_d N_OUT8_Mn9@464_g N_VSS_Mn9@464_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@465 N_OUT9_Mp9@465_d N_OUT8_Mp9@465_g N_VDD_Mp9@465_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@464 N_OUT9_Mp9@464_d N_OUT8_Mp9@464_g N_VDD_Mp9@464_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@463 N_OUT9_Mn9@463_d N_OUT8_Mn9@463_g N_VSS_Mn9@463_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@462 N_OUT9_Mn9@462_d N_OUT8_Mn9@462_g N_VSS_Mn9@462_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@463 N_OUT9_Mp9@463_d N_OUT8_Mp9@463_g N_VDD_Mp9@463_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@462 N_OUT9_Mp9@462_d N_OUT8_Mp9@462_g N_VDD_Mp9@462_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@461 N_OUT9_Mn9@461_d N_OUT8_Mn9@461_g N_VSS_Mn9@461_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@460 N_OUT9_Mn9@460_d N_OUT8_Mn9@460_g N_VSS_Mn9@460_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@461 N_OUT9_Mp9@461_d N_OUT8_Mp9@461_g N_VDD_Mp9@461_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@460 N_OUT9_Mp9@460_d N_OUT8_Mp9@460_g N_VDD_Mp9@460_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@459 N_OUT9_Mn9@459_d N_OUT8_Mn9@459_g N_VSS_Mn9@459_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@458 N_OUT9_Mn9@458_d N_OUT8_Mn9@458_g N_VSS_Mn9@458_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@459 N_OUT9_Mp9@459_d N_OUT8_Mp9@459_g N_VDD_Mp9@459_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@458 N_OUT9_Mp9@458_d N_OUT8_Mp9@458_g N_VDD_Mp9@458_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@457 N_OUT9_Mn9@457_d N_OUT8_Mn9@457_g N_VSS_Mn9@457_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@456 N_OUT9_Mn9@456_d N_OUT8_Mn9@456_g N_VSS_Mn9@456_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@457 N_OUT9_Mp9@457_d N_OUT8_Mp9@457_g N_VDD_Mp9@457_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@456 N_OUT9_Mp9@456_d N_OUT8_Mp9@456_g N_VDD_Mp9@456_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@455 N_OUT9_Mn9@455_d N_OUT8_Mn9@455_g N_VSS_Mn9@455_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@454 N_OUT9_Mn9@454_d N_OUT8_Mn9@454_g N_VSS_Mn9@454_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@455 N_OUT9_Mp9@455_d N_OUT8_Mp9@455_g N_VDD_Mp9@455_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@454 N_OUT9_Mp9@454_d N_OUT8_Mp9@454_g N_VDD_Mp9@454_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@453 N_OUT9_Mn9@453_d N_OUT8_Mn9@453_g N_VSS_Mn9@453_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@452 N_OUT9_Mn9@452_d N_OUT8_Mn9@452_g N_VSS_Mn9@452_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@453 N_OUT9_Mp9@453_d N_OUT8_Mp9@453_g N_VDD_Mp9@453_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@452 N_OUT9_Mp9@452_d N_OUT8_Mp9@452_g N_VDD_Mp9@452_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@451 N_OUT9_Mn9@451_d N_OUT8_Mn9@451_g N_VSS_Mn9@451_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@450 N_OUT9_Mn9@450_d N_OUT8_Mn9@450_g N_VSS_Mn9@450_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@451 N_OUT9_Mp9@451_d N_OUT8_Mp9@451_g N_VDD_Mp9@451_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@450 N_OUT9_Mp9@450_d N_OUT8_Mp9@450_g N_VDD_Mp9@450_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@449 N_OUT9_Mn9@449_d N_OUT8_Mn9@449_g N_VSS_Mn9@449_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@448 N_OUT9_Mn9@448_d N_OUT8_Mn9@448_g N_VSS_Mn9@448_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@449 N_OUT9_Mp9@449_d N_OUT8_Mp9@449_g N_VDD_Mp9@449_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@448 N_OUT9_Mp9@448_d N_OUT8_Mp9@448_g N_VDD_Mp9@448_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@447 N_OUT9_Mn9@447_d N_OUT8_Mn9@447_g N_VSS_Mn9@447_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@446 N_OUT9_Mn9@446_d N_OUT8_Mn9@446_g N_VSS_Mn9@446_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@447 N_OUT9_Mp9@447_d N_OUT8_Mp9@447_g N_VDD_Mp9@447_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@446 N_OUT9_Mp9@446_d N_OUT8_Mp9@446_g N_VDD_Mp9@446_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@445 N_OUT9_Mn9@445_d N_OUT8_Mn9@445_g N_VSS_Mn9@445_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@444 N_OUT9_Mn9@444_d N_OUT8_Mn9@444_g N_VSS_Mn9@444_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@445 N_OUT9_Mp9@445_d N_OUT8_Mp9@445_g N_VDD_Mp9@445_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@444 N_OUT9_Mp9@444_d N_OUT8_Mp9@444_g N_VDD_Mp9@444_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@443 N_OUT9_Mn9@443_d N_OUT8_Mn9@443_g N_VSS_Mn9@443_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@442 N_OUT9_Mn9@442_d N_OUT8_Mn9@442_g N_VSS_Mn9@442_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@443 N_OUT9_Mp9@443_d N_OUT8_Mp9@443_g N_VDD_Mp9@443_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@442 N_OUT9_Mp9@442_d N_OUT8_Mp9@442_g N_VDD_Mp9@442_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@441 N_OUT9_Mn9@441_d N_OUT8_Mn9@441_g N_VSS_Mn9@441_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@440 N_OUT9_Mn9@440_d N_OUT8_Mn9@440_g N_VSS_Mn9@440_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@441 N_OUT9_Mp9@441_d N_OUT8_Mp9@441_g N_VDD_Mp9@441_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@440 N_OUT9_Mp9@440_d N_OUT8_Mp9@440_g N_VDD_Mp9@440_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@439 N_OUT9_Mn9@439_d N_OUT8_Mn9@439_g N_VSS_Mn9@439_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@438 N_OUT9_Mn9@438_d N_OUT8_Mn9@438_g N_VSS_Mn9@438_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@439 N_OUT9_Mp9@439_d N_OUT8_Mp9@439_g N_VDD_Mp9@439_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@438 N_OUT9_Mp9@438_d N_OUT8_Mp9@438_g N_VDD_Mp9@438_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@437 N_OUT9_Mn9@437_d N_OUT8_Mn9@437_g N_VSS_Mn9@437_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@436 N_OUT9_Mn9@436_d N_OUT8_Mn9@436_g N_VSS_Mn9@436_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@437 N_OUT9_Mp9@437_d N_OUT8_Mp9@437_g N_VDD_Mp9@437_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@436 N_OUT9_Mp9@436_d N_OUT8_Mp9@436_g N_VDD_Mp9@436_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@435 N_OUT9_Mn9@435_d N_OUT8_Mn9@435_g N_VSS_Mn9@435_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@434 N_OUT9_Mn9@434_d N_OUT8_Mn9@434_g N_VSS_Mn9@434_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@435 N_OUT9_Mp9@435_d N_OUT8_Mp9@435_g N_VDD_Mp9@435_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@434 N_OUT9_Mp9@434_d N_OUT8_Mp9@434_g N_VDD_Mp9@434_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@433 N_OUT9_Mn9@433_d N_OUT8_Mn9@433_g N_VSS_Mn9@433_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@432 N_OUT9_Mn9@432_d N_OUT8_Mn9@432_g N_VSS_Mn9@432_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@433 N_OUT9_Mp9@433_d N_OUT8_Mp9@433_g N_VDD_Mp9@433_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@432 N_OUT9_Mp9@432_d N_OUT8_Mp9@432_g N_VDD_Mp9@432_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@431 N_OUT9_Mn9@431_d N_OUT8_Mn9@431_g N_VSS_Mn9@431_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@430 N_OUT9_Mn9@430_d N_OUT8_Mn9@430_g N_VSS_Mn9@430_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@431 N_OUT9_Mp9@431_d N_OUT8_Mp9@431_g N_VDD_Mp9@431_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@430 N_OUT9_Mp9@430_d N_OUT8_Mp9@430_g N_VDD_Mp9@430_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@429 N_OUT9_Mn9@429_d N_OUT8_Mn9@429_g N_VSS_Mn9@429_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@428 N_OUT9_Mn9@428_d N_OUT8_Mn9@428_g N_VSS_Mn9@428_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@429 N_OUT9_Mp9@429_d N_OUT8_Mp9@429_g N_VDD_Mp9@429_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@428 N_OUT9_Mp9@428_d N_OUT8_Mp9@428_g N_VDD_Mp9@428_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@427 N_OUT9_Mn9@427_d N_OUT8_Mn9@427_g N_VSS_Mn9@427_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@426 N_OUT9_Mn9@426_d N_OUT8_Mn9@426_g N_VSS_Mn9@426_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@427 N_OUT9_Mp9@427_d N_OUT8_Mp9@427_g N_VDD_Mp9@427_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@426 N_OUT9_Mp9@426_d N_OUT8_Mp9@426_g N_VDD_Mp9@426_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@425 N_OUT9_Mn9@425_d N_OUT8_Mn9@425_g N_VSS_Mn9@425_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@424 N_OUT9_Mn9@424_d N_OUT8_Mn9@424_g N_VSS_Mn9@424_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@425 N_OUT9_Mp9@425_d N_OUT8_Mp9@425_g N_VDD_Mp9@425_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@424 N_OUT9_Mp9@424_d N_OUT8_Mp9@424_g N_VDD_Mp9@424_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@423 N_OUT9_Mn9@423_d N_OUT8_Mn9@423_g N_VSS_Mn9@423_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@422 N_OUT9_Mn9@422_d N_OUT8_Mn9@422_g N_VSS_Mn9@422_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@423 N_OUT9_Mp9@423_d N_OUT8_Mp9@423_g N_VDD_Mp9@423_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@422 N_OUT9_Mp9@422_d N_OUT8_Mp9@422_g N_VDD_Mp9@422_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@421 N_OUT9_Mn9@421_d N_OUT8_Mn9@421_g N_VSS_Mn9@421_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@420 N_OUT9_Mn9@420_d N_OUT8_Mn9@420_g N_VSS_Mn9@420_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@421 N_OUT9_Mp9@421_d N_OUT8_Mp9@421_g N_VDD_Mp9@421_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@420 N_OUT9_Mp9@420_d N_OUT8_Mp9@420_g N_VDD_Mp9@420_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@419 N_OUT9_Mn9@419_d N_OUT8_Mn9@419_g N_VSS_Mn9@419_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@418 N_OUT9_Mn9@418_d N_OUT8_Mn9@418_g N_VSS_Mn9@418_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@419 N_OUT9_Mp9@419_d N_OUT8_Mp9@419_g N_VDD_Mp9@419_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@418 N_OUT9_Mp9@418_d N_OUT8_Mp9@418_g N_VDD_Mp9@418_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@417 N_OUT9_Mn9@417_d N_OUT8_Mn9@417_g N_VSS_Mn9@417_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@416 N_OUT9_Mn9@416_d N_OUT8_Mn9@416_g N_VSS_Mn9@416_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@417 N_OUT9_Mp9@417_d N_OUT8_Mp9@417_g N_VDD_Mp9@417_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@416 N_OUT9_Mp9@416_d N_OUT8_Mp9@416_g N_VDD_Mp9@416_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@415 N_OUT9_Mn9@415_d N_OUT8_Mn9@415_g N_VSS_Mn9@415_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@414 N_OUT9_Mn9@414_d N_OUT8_Mn9@414_g N_VSS_Mn9@414_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@415 N_OUT9_Mp9@415_d N_OUT8_Mp9@415_g N_VDD_Mp9@415_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@414 N_OUT9_Mp9@414_d N_OUT8_Mp9@414_g N_VDD_Mp9@414_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@413 N_OUT9_Mn9@413_d N_OUT8_Mn9@413_g N_VSS_Mn9@413_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@412 N_OUT9_Mn9@412_d N_OUT8_Mn9@412_g N_VSS_Mn9@412_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@413 N_OUT9_Mp9@413_d N_OUT8_Mp9@413_g N_VDD_Mp9@413_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@412 N_OUT9_Mp9@412_d N_OUT8_Mp9@412_g N_VDD_Mp9@412_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@411 N_OUT9_Mn9@411_d N_OUT8_Mn9@411_g N_VSS_Mn9@411_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@410 N_OUT9_Mn9@410_d N_OUT8_Mn9@410_g N_VSS_Mn9@410_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@411 N_OUT9_Mp9@411_d N_OUT8_Mp9@411_g N_VDD_Mp9@411_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@410 N_OUT9_Mp9@410_d N_OUT8_Mp9@410_g N_VDD_Mp9@410_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@409 N_OUT9_Mn9@409_d N_OUT8_Mn9@409_g N_VSS_Mn9@409_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@408 N_OUT9_Mn9@408_d N_OUT8_Mn9@408_g N_VSS_Mn9@408_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@409 N_OUT9_Mp9@409_d N_OUT8_Mp9@409_g N_VDD_Mp9@409_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@408 N_OUT9_Mp9@408_d N_OUT8_Mp9@408_g N_VDD_Mp9@408_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@407 N_OUT9_Mn9@407_d N_OUT8_Mn9@407_g N_VSS_Mn9@407_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@406 N_OUT9_Mn9@406_d N_OUT8_Mn9@406_g N_VSS_Mn9@406_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@407 N_OUT9_Mp9@407_d N_OUT8_Mp9@407_g N_VDD_Mp9@407_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@406 N_OUT9_Mp9@406_d N_OUT8_Mp9@406_g N_VDD_Mp9@406_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@405 N_OUT9_Mn9@405_d N_OUT8_Mn9@405_g N_VSS_Mn9@405_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@404 N_OUT9_Mn9@404_d N_OUT8_Mn9@404_g N_VSS_Mn9@404_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@405 N_OUT9_Mp9@405_d N_OUT8_Mp9@405_g N_VDD_Mp9@405_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@404 N_OUT9_Mp9@404_d N_OUT8_Mp9@404_g N_VDD_Mp9@404_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@403 N_OUT9_Mn9@403_d N_OUT8_Mn9@403_g N_VSS_Mn9@403_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@402 N_OUT9_Mn9@402_d N_OUT8_Mn9@402_g N_VSS_Mn9@402_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@403 N_OUT9_Mp9@403_d N_OUT8_Mp9@403_g N_VDD_Mp9@403_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@402 N_OUT9_Mp9@402_d N_OUT8_Mp9@402_g N_VDD_Mp9@402_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@401 N_OUT9_Mn9@401_d N_OUT8_Mn9@401_g N_VSS_Mn9@401_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@400 N_OUT9_Mn9@400_d N_OUT8_Mn9@400_g N_VSS_Mn9@400_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@401 N_OUT9_Mp9@401_d N_OUT8_Mp9@401_g N_VDD_Mp9@401_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@400 N_OUT9_Mp9@400_d N_OUT8_Mp9@400_g N_VDD_Mp9@400_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@399 N_OUT9_Mn9@399_d N_OUT8_Mn9@399_g N_VSS_Mn9@399_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@398 N_OUT9_Mn9@398_d N_OUT8_Mn9@398_g N_VSS_Mn9@398_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@399 N_OUT9_Mp9@399_d N_OUT8_Mp9@399_g N_VDD_Mp9@399_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@398 N_OUT9_Mp9@398_d N_OUT8_Mp9@398_g N_VDD_Mp9@398_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@397 N_OUT9_Mn9@397_d N_OUT8_Mn9@397_g N_VSS_Mn9@397_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@396 N_OUT9_Mn9@396_d N_OUT8_Mn9@396_g N_VSS_Mn9@396_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@397 N_OUT9_Mp9@397_d N_OUT8_Mp9@397_g N_VDD_Mp9@397_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@396 N_OUT9_Mp9@396_d N_OUT8_Mp9@396_g N_VDD_Mp9@396_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@395 N_OUT9_Mn9@395_d N_OUT8_Mn9@395_g N_VSS_Mn9@395_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@394 N_OUT9_Mn9@394_d N_OUT8_Mn9@394_g N_VSS_Mn9@394_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@395 N_OUT9_Mp9@395_d N_OUT8_Mp9@395_g N_VDD_Mp9@395_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@394 N_OUT9_Mp9@394_d N_OUT8_Mp9@394_g N_VDD_Mp9@394_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@393 N_OUT9_Mn9@393_d N_OUT8_Mn9@393_g N_VSS_Mn9@393_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@392 N_OUT9_Mn9@392_d N_OUT8_Mn9@392_g N_VSS_Mn9@392_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@393 N_OUT9_Mp9@393_d N_OUT8_Mp9@393_g N_VDD_Mp9@393_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@392 N_OUT9_Mp9@392_d N_OUT8_Mp9@392_g N_VDD_Mp9@392_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@391 N_OUT9_Mn9@391_d N_OUT8_Mn9@391_g N_VSS_Mn9@391_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@390 N_OUT9_Mn9@390_d N_OUT8_Mn9@390_g N_VSS_Mn9@390_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@391 N_OUT9_Mp9@391_d N_OUT8_Mp9@391_g N_VDD_Mp9@391_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@390 N_OUT9_Mp9@390_d N_OUT8_Mp9@390_g N_VDD_Mp9@390_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@389 N_OUT9_Mn9@389_d N_OUT8_Mn9@389_g N_VSS_Mn9@389_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@388 N_OUT9_Mn9@388_d N_OUT8_Mn9@388_g N_VSS_Mn9@388_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@389 N_OUT9_Mp9@389_d N_OUT8_Mp9@389_g N_VDD_Mp9@389_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@388 N_OUT9_Mp9@388_d N_OUT8_Mp9@388_g N_VDD_Mp9@388_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@387 N_OUT9_Mn9@387_d N_OUT8_Mn9@387_g N_VSS_Mn9@387_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@386 N_OUT9_Mn9@386_d N_OUT8_Mn9@386_g N_VSS_Mn9@386_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@387 N_OUT9_Mp9@387_d N_OUT8_Mp9@387_g N_VDD_Mp9@387_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@386 N_OUT9_Mp9@386_d N_OUT8_Mp9@386_g N_VDD_Mp9@386_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@385 N_OUT9_Mn9@385_d N_OUT8_Mn9@385_g N_VSS_Mn9@385_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@384 N_OUT9_Mn9@384_d N_OUT8_Mn9@384_g N_VSS_Mn9@384_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@385 N_OUT9_Mp9@385_d N_OUT8_Mp9@385_g N_VDD_Mp9@385_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@384 N_OUT9_Mp9@384_d N_OUT8_Mp9@384_g N_VDD_Mp9@384_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@383 N_OUT9_Mn9@383_d N_OUT8_Mn9@383_g N_VSS_Mn9@383_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@382 N_OUT9_Mn9@382_d N_OUT8_Mn9@382_g N_VSS_Mn9@382_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@383 N_OUT9_Mp9@383_d N_OUT8_Mp9@383_g N_VDD_Mp9@383_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@382 N_OUT9_Mp9@382_d N_OUT8_Mp9@382_g N_VDD_Mp9@382_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@381 N_OUT9_Mn9@381_d N_OUT8_Mn9@381_g N_VSS_Mn9@381_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@380 N_OUT9_Mn9@380_d N_OUT8_Mn9@380_g N_VSS_Mn9@380_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@381 N_OUT9_Mp9@381_d N_OUT8_Mp9@381_g N_VDD_Mp9@381_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@380 N_OUT9_Mp9@380_d N_OUT8_Mp9@380_g N_VDD_Mp9@380_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@379 N_OUT9_Mn9@379_d N_OUT8_Mn9@379_g N_VSS_Mn9@379_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@378 N_OUT9_Mn9@378_d N_OUT8_Mn9@378_g N_VSS_Mn9@378_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@379 N_OUT9_Mp9@379_d N_OUT8_Mp9@379_g N_VDD_Mp9@379_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@378 N_OUT9_Mp9@378_d N_OUT8_Mp9@378_g N_VDD_Mp9@378_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@377 N_OUT9_Mn9@377_d N_OUT8_Mn9@377_g N_VSS_Mn9@377_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@376 N_OUT9_Mn9@376_d N_OUT8_Mn9@376_g N_VSS_Mn9@376_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@377 N_OUT9_Mp9@377_d N_OUT8_Mp9@377_g N_VDD_Mp9@377_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@376 N_OUT9_Mp9@376_d N_OUT8_Mp9@376_g N_VDD_Mp9@376_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@375 N_OUT9_Mn9@375_d N_OUT8_Mn9@375_g N_VSS_Mn9@375_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@374 N_OUT9_Mn9@374_d N_OUT8_Mn9@374_g N_VSS_Mn9@374_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@375 N_OUT9_Mp9@375_d N_OUT8_Mp9@375_g N_VDD_Mp9@375_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@374 N_OUT9_Mp9@374_d N_OUT8_Mp9@374_g N_VDD_Mp9@374_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@373 N_OUT9_Mn9@373_d N_OUT8_Mn9@373_g N_VSS_Mn9@373_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@372 N_OUT9_Mn9@372_d N_OUT8_Mn9@372_g N_VSS_Mn9@372_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@373 N_OUT9_Mp9@373_d N_OUT8_Mp9@373_g N_VDD_Mp9@373_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@372 N_OUT9_Mp9@372_d N_OUT8_Mp9@372_g N_VDD_Mp9@372_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@371 N_OUT9_Mn9@371_d N_OUT8_Mn9@371_g N_VSS_Mn9@371_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@370 N_OUT9_Mn9@370_d N_OUT8_Mn9@370_g N_VSS_Mn9@370_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@371 N_OUT9_Mp9@371_d N_OUT8_Mp9@371_g N_VDD_Mp9@371_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@370 N_OUT9_Mp9@370_d N_OUT8_Mp9@370_g N_VDD_Mp9@370_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@369 N_OUT9_Mn9@369_d N_OUT8_Mn9@369_g N_VSS_Mn9@369_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@368 N_OUT9_Mn9@368_d N_OUT8_Mn9@368_g N_VSS_Mn9@368_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@369 N_OUT9_Mp9@369_d N_OUT8_Mp9@369_g N_VDD_Mp9@369_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@368 N_OUT9_Mp9@368_d N_OUT8_Mp9@368_g N_VDD_Mp9@368_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@367 N_OUT9_Mn9@367_d N_OUT8_Mn9@367_g N_VSS_Mn9@367_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@366 N_OUT9_Mn9@366_d N_OUT8_Mn9@366_g N_VSS_Mn9@366_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@367 N_OUT9_Mp9@367_d N_OUT8_Mp9@367_g N_VDD_Mp9@367_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@366 N_OUT9_Mp9@366_d N_OUT8_Mp9@366_g N_VDD_Mp9@366_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@365 N_OUT9_Mn9@365_d N_OUT8_Mn9@365_g N_VSS_Mn9@365_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@364 N_OUT9_Mn9@364_d N_OUT8_Mn9@364_g N_VSS_Mn9@364_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@365 N_OUT9_Mp9@365_d N_OUT8_Mp9@365_g N_VDD_Mp9@365_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@364 N_OUT9_Mp9@364_d N_OUT8_Mp9@364_g N_VDD_Mp9@364_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@363 N_OUT9_Mn9@363_d N_OUT8_Mn9@363_g N_VSS_Mn9@363_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@362 N_OUT9_Mn9@362_d N_OUT8_Mn9@362_g N_VSS_Mn9@362_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@363 N_OUT9_Mp9@363_d N_OUT8_Mp9@363_g N_VDD_Mp9@363_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@362 N_OUT9_Mp9@362_d N_OUT8_Mp9@362_g N_VDD_Mp9@362_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@361 N_OUT9_Mn9@361_d N_OUT8_Mn9@361_g N_VSS_Mn9@361_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@360 N_OUT9_Mn9@360_d N_OUT8_Mn9@360_g N_VSS_Mn9@360_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@361 N_OUT9_Mp9@361_d N_OUT8_Mp9@361_g N_VDD_Mp9@361_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@360 N_OUT9_Mp9@360_d N_OUT8_Mp9@360_g N_VDD_Mp9@360_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@359 N_OUT9_Mn9@359_d N_OUT8_Mn9@359_g N_VSS_Mn9@359_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@358 N_OUT9_Mn9@358_d N_OUT8_Mn9@358_g N_VSS_Mn9@358_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@359 N_OUT9_Mp9@359_d N_OUT8_Mp9@359_g N_VDD_Mp9@359_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@358 N_OUT9_Mp9@358_d N_OUT8_Mp9@358_g N_VDD_Mp9@358_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@357 N_OUT9_Mn9@357_d N_OUT8_Mn9@357_g N_VSS_Mn9@357_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@356 N_OUT9_Mn9@356_d N_OUT8_Mn9@356_g N_VSS_Mn9@356_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@357 N_OUT9_Mp9@357_d N_OUT8_Mp9@357_g N_VDD_Mp9@357_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@356 N_OUT9_Mp9@356_d N_OUT8_Mp9@356_g N_VDD_Mp9@356_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@355 N_OUT9_Mn9@355_d N_OUT8_Mn9@355_g N_VSS_Mn9@355_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@354 N_OUT9_Mn9@354_d N_OUT8_Mn9@354_g N_VSS_Mn9@354_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@355 N_OUT9_Mp9@355_d N_OUT8_Mp9@355_g N_VDD_Mp9@355_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@354 N_OUT9_Mp9@354_d N_OUT8_Mp9@354_g N_VDD_Mp9@354_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@353 N_OUT9_Mn9@353_d N_OUT8_Mn9@353_g N_VSS_Mn9@353_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@352 N_OUT9_Mn9@352_d N_OUT8_Mn9@352_g N_VSS_Mn9@352_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@353 N_OUT9_Mp9@353_d N_OUT8_Mp9@353_g N_VDD_Mp9@353_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@352 N_OUT9_Mp9@352_d N_OUT8_Mp9@352_g N_VDD_Mp9@352_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@351 N_OUT9_Mn9@351_d N_OUT8_Mn9@351_g N_VSS_Mn9@351_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@350 N_OUT9_Mn9@350_d N_OUT8_Mn9@350_g N_VSS_Mn9@350_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@351 N_OUT9_Mp9@351_d N_OUT8_Mp9@351_g N_VDD_Mp9@351_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@350 N_OUT9_Mp9@350_d N_OUT8_Mp9@350_g N_VDD_Mp9@350_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@349 N_OUT9_Mn9@349_d N_OUT8_Mn9@349_g N_VSS_Mn9@349_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@348 N_OUT9_Mn9@348_d N_OUT8_Mn9@348_g N_VSS_Mn9@348_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@349 N_OUT9_Mp9@349_d N_OUT8_Mp9@349_g N_VDD_Mp9@349_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@348 N_OUT9_Mp9@348_d N_OUT8_Mp9@348_g N_VDD_Mp9@348_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@347 N_OUT9_Mn9@347_d N_OUT8_Mn9@347_g N_VSS_Mn9@347_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@346 N_OUT9_Mn9@346_d N_OUT8_Mn9@346_g N_VSS_Mn9@346_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@347 N_OUT9_Mp9@347_d N_OUT8_Mp9@347_g N_VDD_Mp9@347_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@346 N_OUT9_Mp9@346_d N_OUT8_Mp9@346_g N_VDD_Mp9@346_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@345 N_OUT9_Mn9@345_d N_OUT8_Mn9@345_g N_VSS_Mn9@345_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@344 N_OUT9_Mn9@344_d N_OUT8_Mn9@344_g N_VSS_Mn9@344_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@345 N_OUT9_Mp9@345_d N_OUT8_Mp9@345_g N_VDD_Mp9@345_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@344 N_OUT9_Mp9@344_d N_OUT8_Mp9@344_g N_VDD_Mp9@344_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@343 N_OUT9_Mn9@343_d N_OUT8_Mn9@343_g N_VSS_Mn9@343_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@342 N_OUT9_Mn9@342_d N_OUT8_Mn9@342_g N_VSS_Mn9@342_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@343 N_OUT9_Mp9@343_d N_OUT8_Mp9@343_g N_VDD_Mp9@343_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@342 N_OUT9_Mp9@342_d N_OUT8_Mp9@342_g N_VDD_Mp9@342_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@341 N_OUT9_Mn9@341_d N_OUT8_Mn9@341_g N_VSS_Mn9@341_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@340 N_OUT9_Mn9@340_d N_OUT8_Mn9@340_g N_VSS_Mn9@340_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@341 N_OUT9_Mp9@341_d N_OUT8_Mp9@341_g N_VDD_Mp9@341_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@340 N_OUT9_Mp9@340_d N_OUT8_Mp9@340_g N_VDD_Mp9@340_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@339 N_OUT9_Mn9@339_d N_OUT8_Mn9@339_g N_VSS_Mn9@339_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@338 N_OUT9_Mn9@338_d N_OUT8_Mn9@338_g N_VSS_Mn9@338_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@339 N_OUT9_Mp9@339_d N_OUT8_Mp9@339_g N_VDD_Mp9@339_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@338 N_OUT9_Mp9@338_d N_OUT8_Mp9@338_g N_VDD_Mp9@338_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@337 N_OUT9_Mn9@337_d N_OUT8_Mn9@337_g N_VSS_Mn9@337_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@336 N_OUT9_Mn9@336_d N_OUT8_Mn9@336_g N_VSS_Mn9@336_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@337 N_OUT9_Mp9@337_d N_OUT8_Mp9@337_g N_VDD_Mp9@337_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@336 N_OUT9_Mp9@336_d N_OUT8_Mp9@336_g N_VDD_Mp9@336_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@335 N_OUT9_Mn9@335_d N_OUT8_Mn9@335_g N_VSS_Mn9@335_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@334 N_OUT9_Mn9@334_d N_OUT8_Mn9@334_g N_VSS_Mn9@334_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@335 N_OUT9_Mp9@335_d N_OUT8_Mp9@335_g N_VDD_Mp9@335_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@334 N_OUT9_Mp9@334_d N_OUT8_Mp9@334_g N_VDD_Mp9@334_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@333 N_OUT9_Mn9@333_d N_OUT8_Mn9@333_g N_VSS_Mn9@333_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@332 N_OUT9_Mn9@332_d N_OUT8_Mn9@332_g N_VSS_Mn9@332_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@333 N_OUT9_Mp9@333_d N_OUT8_Mp9@333_g N_VDD_Mp9@333_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@332 N_OUT9_Mp9@332_d N_OUT8_Mp9@332_g N_VDD_Mp9@332_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@331 N_OUT9_Mn9@331_d N_OUT8_Mn9@331_g N_VSS_Mn9@331_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@330 N_OUT9_Mn9@330_d N_OUT8_Mn9@330_g N_VSS_Mn9@330_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@331 N_OUT9_Mp9@331_d N_OUT8_Mp9@331_g N_VDD_Mp9@331_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@330 N_OUT9_Mp9@330_d N_OUT8_Mp9@330_g N_VDD_Mp9@330_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@329 N_OUT9_Mn9@329_d N_OUT8_Mn9@329_g N_VSS_Mn9@329_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@328 N_OUT9_Mn9@328_d N_OUT8_Mn9@328_g N_VSS_Mn9@328_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@329 N_OUT9_Mp9@329_d N_OUT8_Mp9@329_g N_VDD_Mp9@329_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@328 N_OUT9_Mp9@328_d N_OUT8_Mp9@328_g N_VDD_Mp9@328_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@327 N_OUT9_Mn9@327_d N_OUT8_Mn9@327_g N_VSS_Mn9@327_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@326 N_OUT9_Mn9@326_d N_OUT8_Mn9@326_g N_VSS_Mn9@326_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@327 N_OUT9_Mp9@327_d N_OUT8_Mp9@327_g N_VDD_Mp9@327_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@326 N_OUT9_Mp9@326_d N_OUT8_Mp9@326_g N_VDD_Mp9@326_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@325 N_OUT9_Mn9@325_d N_OUT8_Mn9@325_g N_VSS_Mn9@325_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@324 N_OUT9_Mn9@324_d N_OUT8_Mn9@324_g N_VSS_Mn9@324_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@325 N_OUT9_Mp9@325_d N_OUT8_Mp9@325_g N_VDD_Mp9@325_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@324 N_OUT9_Mp9@324_d N_OUT8_Mp9@324_g N_VDD_Mp9@324_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@323 N_OUT9_Mn9@323_d N_OUT8_Mn9@323_g N_VSS_Mn9@323_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@322 N_OUT9_Mn9@322_d N_OUT8_Mn9@322_g N_VSS_Mn9@322_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@323 N_OUT9_Mp9@323_d N_OUT8_Mp9@323_g N_VDD_Mp9@323_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@322 N_OUT9_Mp9@322_d N_OUT8_Mp9@322_g N_VDD_Mp9@322_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@321 N_OUT9_Mn9@321_d N_OUT8_Mn9@321_g N_VSS_Mn9@321_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@320 N_OUT9_Mn9@320_d N_OUT8_Mn9@320_g N_VSS_Mn9@320_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@321 N_OUT9_Mp9@321_d N_OUT8_Mp9@321_g N_VDD_Mp9@321_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@320 N_OUT9_Mp9@320_d N_OUT8_Mp9@320_g N_VDD_Mp9@320_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@319 N_OUT9_Mn9@319_d N_OUT8_Mn9@319_g N_VSS_Mn9@319_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@318 N_OUT9_Mn9@318_d N_OUT8_Mn9@318_g N_VSS_Mn9@318_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@319 N_OUT9_Mp9@319_d N_OUT8_Mp9@319_g N_VDD_Mp9@319_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@318 N_OUT9_Mp9@318_d N_OUT8_Mp9@318_g N_VDD_Mp9@318_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@317 N_OUT9_Mn9@317_d N_OUT8_Mn9@317_g N_VSS_Mn9@317_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@316 N_OUT9_Mn9@316_d N_OUT8_Mn9@316_g N_VSS_Mn9@316_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@317 N_OUT9_Mp9@317_d N_OUT8_Mp9@317_g N_VDD_Mp9@317_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@316 N_OUT9_Mp9@316_d N_OUT8_Mp9@316_g N_VDD_Mp9@316_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@315 N_OUT9_Mn9@315_d N_OUT8_Mn9@315_g N_VSS_Mn9@315_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@314 N_OUT9_Mn9@314_d N_OUT8_Mn9@314_g N_VSS_Mn9@314_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@315 N_OUT9_Mp9@315_d N_OUT8_Mp9@315_g N_VDD_Mp9@315_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@314 N_OUT9_Mp9@314_d N_OUT8_Mp9@314_g N_VDD_Mp9@314_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@313 N_OUT9_Mn9@313_d N_OUT8_Mn9@313_g N_VSS_Mn9@313_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@312 N_OUT9_Mn9@312_d N_OUT8_Mn9@312_g N_VSS_Mn9@312_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@313 N_OUT9_Mp9@313_d N_OUT8_Mp9@313_g N_VDD_Mp9@313_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@312 N_OUT9_Mp9@312_d N_OUT8_Mp9@312_g N_VDD_Mp9@312_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@311 N_OUT9_Mn9@311_d N_OUT8_Mn9@311_g N_VSS_Mn9@311_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@310 N_OUT9_Mn9@310_d N_OUT8_Mn9@310_g N_VSS_Mn9@310_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@311 N_OUT9_Mp9@311_d N_OUT8_Mp9@311_g N_VDD_Mp9@311_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@310 N_OUT9_Mp9@310_d N_OUT8_Mp9@310_g N_VDD_Mp9@310_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@309 N_OUT9_Mn9@309_d N_OUT8_Mn9@309_g N_VSS_Mn9@309_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@308 N_OUT9_Mn9@308_d N_OUT8_Mn9@308_g N_VSS_Mn9@308_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@309 N_OUT9_Mp9@309_d N_OUT8_Mp9@309_g N_VDD_Mp9@309_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@308 N_OUT9_Mp9@308_d N_OUT8_Mp9@308_g N_VDD_Mp9@308_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@307 N_OUT9_Mn9@307_d N_OUT8_Mn9@307_g N_VSS_Mn9@307_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@306 N_OUT9_Mn9@306_d N_OUT8_Mn9@306_g N_VSS_Mn9@306_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@307 N_OUT9_Mp9@307_d N_OUT8_Mp9@307_g N_VDD_Mp9@307_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@306 N_OUT9_Mp9@306_d N_OUT8_Mp9@306_g N_VDD_Mp9@306_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@305 N_OUT9_Mn9@305_d N_OUT8_Mn9@305_g N_VSS_Mn9@305_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@304 N_OUT9_Mn9@304_d N_OUT8_Mn9@304_g N_VSS_Mn9@304_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@305 N_OUT9_Mp9@305_d N_OUT8_Mp9@305_g N_VDD_Mp9@305_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@304 N_OUT9_Mp9@304_d N_OUT8_Mp9@304_g N_VDD_Mp9@304_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@303 N_OUT9_Mn9@303_d N_OUT8_Mn9@303_g N_VSS_Mn9@303_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@302 N_OUT9_Mn9@302_d N_OUT8_Mn9@302_g N_VSS_Mn9@302_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@303 N_OUT9_Mp9@303_d N_OUT8_Mp9@303_g N_VDD_Mp9@303_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@302 N_OUT9_Mp9@302_d N_OUT8_Mp9@302_g N_VDD_Mp9@302_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@301 N_OUT9_Mn9@301_d N_OUT8_Mn9@301_g N_VSS_Mn9@301_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@300 N_OUT9_Mn9@300_d N_OUT8_Mn9@300_g N_VSS_Mn9@300_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@301 N_OUT9_Mp9@301_d N_OUT8_Mp9@301_g N_VDD_Mp9@301_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@300 N_OUT9_Mp9@300_d N_OUT8_Mp9@300_g N_VDD_Mp9@300_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@299 N_OUT9_Mn9@299_d N_OUT8_Mn9@299_g N_VSS_Mn9@299_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@298 N_OUT9_Mn9@298_d N_OUT8_Mn9@298_g N_VSS_Mn9@298_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@299 N_OUT9_Mp9@299_d N_OUT8_Mp9@299_g N_VDD_Mp9@299_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@298 N_OUT9_Mp9@298_d N_OUT8_Mp9@298_g N_VDD_Mp9@298_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@297 N_OUT9_Mn9@297_d N_OUT8_Mn9@297_g N_VSS_Mn9@297_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@296 N_OUT9_Mn9@296_d N_OUT8_Mn9@296_g N_VSS_Mn9@296_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@297 N_OUT9_Mp9@297_d N_OUT8_Mp9@297_g N_VDD_Mp9@297_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@296 N_OUT9_Mp9@296_d N_OUT8_Mp9@296_g N_VDD_Mp9@296_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@295 N_OUT9_Mn9@295_d N_OUT8_Mn9@295_g N_VSS_Mn9@295_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@294 N_OUT9_Mn9@294_d N_OUT8_Mn9@294_g N_VSS_Mn9@294_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@295 N_OUT9_Mp9@295_d N_OUT8_Mp9@295_g N_VDD_Mp9@295_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@294 N_OUT9_Mp9@294_d N_OUT8_Mp9@294_g N_VDD_Mp9@294_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@293 N_OUT9_Mn9@293_d N_OUT8_Mn9@293_g N_VSS_Mn9@293_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@292 N_OUT9_Mn9@292_d N_OUT8_Mn9@292_g N_VSS_Mn9@292_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@293 N_OUT9_Mp9@293_d N_OUT8_Mp9@293_g N_VDD_Mp9@293_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@292 N_OUT9_Mp9@292_d N_OUT8_Mp9@292_g N_VDD_Mp9@292_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@291 N_OUT9_Mn9@291_d N_OUT8_Mn9@291_g N_VSS_Mn9@291_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@290 N_OUT9_Mn9@290_d N_OUT8_Mn9@290_g N_VSS_Mn9@290_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@291 N_OUT9_Mp9@291_d N_OUT8_Mp9@291_g N_VDD_Mp9@291_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@290 N_OUT9_Mp9@290_d N_OUT8_Mp9@290_g N_VDD_Mp9@290_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@289 N_OUT9_Mn9@289_d N_OUT8_Mn9@289_g N_VSS_Mn9@289_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@288 N_OUT9_Mn9@288_d N_OUT8_Mn9@288_g N_VSS_Mn9@288_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@289 N_OUT9_Mp9@289_d N_OUT8_Mp9@289_g N_VDD_Mp9@289_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@288 N_OUT9_Mp9@288_d N_OUT8_Mp9@288_g N_VDD_Mp9@288_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@287 N_OUT9_Mn9@287_d N_OUT8_Mn9@287_g N_VSS_Mn9@287_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@286 N_OUT9_Mn9@286_d N_OUT8_Mn9@286_g N_VSS_Mn9@286_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@287 N_OUT9_Mp9@287_d N_OUT8_Mp9@287_g N_VDD_Mp9@287_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@286 N_OUT9_Mp9@286_d N_OUT8_Mp9@286_g N_VDD_Mp9@286_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@285 N_OUT9_Mn9@285_d N_OUT8_Mn9@285_g N_VSS_Mn9@285_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@284 N_OUT9_Mn9@284_d N_OUT8_Mn9@284_g N_VSS_Mn9@284_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@285 N_OUT9_Mp9@285_d N_OUT8_Mp9@285_g N_VDD_Mp9@285_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@284 N_OUT9_Mp9@284_d N_OUT8_Mp9@284_g N_VDD_Mp9@284_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@283 N_OUT9_Mn9@283_d N_OUT8_Mn9@283_g N_VSS_Mn9@283_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@282 N_OUT9_Mn9@282_d N_OUT8_Mn9@282_g N_VSS_Mn9@282_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@283 N_OUT9_Mp9@283_d N_OUT8_Mp9@283_g N_VDD_Mp9@283_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@282 N_OUT9_Mp9@282_d N_OUT8_Mp9@282_g N_VDD_Mp9@282_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@281 N_OUT9_Mn9@281_d N_OUT8_Mn9@281_g N_VSS_Mn9@281_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@280 N_OUT9_Mn9@280_d N_OUT8_Mn9@280_g N_VSS_Mn9@280_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@281 N_OUT9_Mp9@281_d N_OUT8_Mp9@281_g N_VDD_Mp9@281_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@280 N_OUT9_Mp9@280_d N_OUT8_Mp9@280_g N_VDD_Mp9@280_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@279 N_OUT9_Mn9@279_d N_OUT8_Mn9@279_g N_VSS_Mn9@279_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@278 N_OUT9_Mn9@278_d N_OUT8_Mn9@278_g N_VSS_Mn9@278_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@279 N_OUT9_Mp9@279_d N_OUT8_Mp9@279_g N_VDD_Mp9@279_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@278 N_OUT9_Mp9@278_d N_OUT8_Mp9@278_g N_VDD_Mp9@278_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@277 N_OUT9_Mn9@277_d N_OUT8_Mn9@277_g N_VSS_Mn9@277_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@276 N_OUT9_Mn9@276_d N_OUT8_Mn9@276_g N_VSS_Mn9@276_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@277 N_OUT9_Mp9@277_d N_OUT8_Mp9@277_g N_VDD_Mp9@277_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@276 N_OUT9_Mp9@276_d N_OUT8_Mp9@276_g N_VDD_Mp9@276_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@275 N_OUT9_Mn9@275_d N_OUT8_Mn9@275_g N_VSS_Mn9@275_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@274 N_OUT9_Mn9@274_d N_OUT8_Mn9@274_g N_VSS_Mn9@274_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@275 N_OUT9_Mp9@275_d N_OUT8_Mp9@275_g N_VDD_Mp9@275_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@274 N_OUT9_Mp9@274_d N_OUT8_Mp9@274_g N_VDD_Mp9@274_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@273 N_OUT9_Mn9@273_d N_OUT8_Mn9@273_g N_VSS_Mn9@273_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@272 N_OUT9_Mn9@272_d N_OUT8_Mn9@272_g N_VSS_Mn9@272_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@273 N_OUT9_Mp9@273_d N_OUT8_Mp9@273_g N_VDD_Mp9@273_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@272 N_OUT9_Mp9@272_d N_OUT8_Mp9@272_g N_VDD_Mp9@272_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@271 N_OUT9_Mn9@271_d N_OUT8_Mn9@271_g N_VSS_Mn9@271_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@270 N_OUT9_Mn9@270_d N_OUT8_Mn9@270_g N_VSS_Mn9@270_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@271 N_OUT9_Mp9@271_d N_OUT8_Mp9@271_g N_VDD_Mp9@271_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@270 N_OUT9_Mp9@270_d N_OUT8_Mp9@270_g N_VDD_Mp9@270_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@269 N_OUT9_Mn9@269_d N_OUT8_Mn9@269_g N_VSS_Mn9@269_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@268 N_OUT9_Mn9@268_d N_OUT8_Mn9@268_g N_VSS_Mn9@268_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@269 N_OUT9_Mp9@269_d N_OUT8_Mp9@269_g N_VDD_Mp9@269_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@268 N_OUT9_Mp9@268_d N_OUT8_Mp9@268_g N_VDD_Mp9@268_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@267 N_OUT9_Mn9@267_d N_OUT8_Mn9@267_g N_VSS_Mn9@267_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@266 N_OUT9_Mn9@266_d N_OUT8_Mn9@266_g N_VSS_Mn9@266_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@267 N_OUT9_Mp9@267_d N_OUT8_Mp9@267_g N_VDD_Mp9@267_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@266 N_OUT9_Mp9@266_d N_OUT8_Mp9@266_g N_VDD_Mp9@266_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@265 N_OUT9_Mn9@265_d N_OUT8_Mn9@265_g N_VSS_Mn9@265_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@264 N_OUT9_Mn9@264_d N_OUT8_Mn9@264_g N_VSS_Mn9@264_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@265 N_OUT9_Mp9@265_d N_OUT8_Mp9@265_g N_VDD_Mp9@265_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@264 N_OUT9_Mp9@264_d N_OUT8_Mp9@264_g N_VDD_Mp9@264_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@263 N_OUT9_Mn9@263_d N_OUT8_Mn9@263_g N_VSS_Mn9@263_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@262 N_OUT9_Mn9@262_d N_OUT8_Mn9@262_g N_VSS_Mn9@262_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@263 N_OUT9_Mp9@263_d N_OUT8_Mp9@263_g N_VDD_Mp9@263_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@262 N_OUT9_Mp9@262_d N_OUT8_Mp9@262_g N_VDD_Mp9@262_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@261 N_OUT9_Mn9@261_d N_OUT8_Mn9@261_g N_VSS_Mn9@261_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@260 N_OUT9_Mn9@260_d N_OUT8_Mn9@260_g N_VSS_Mn9@260_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@261 N_OUT9_Mp9@261_d N_OUT8_Mp9@261_g N_VDD_Mp9@261_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@260 N_OUT9_Mp9@260_d N_OUT8_Mp9@260_g N_VDD_Mp9@260_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@259 N_OUT9_Mn9@259_d N_OUT8_Mn9@259_g N_VSS_Mn9@259_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@258 N_OUT9_Mn9@258_d N_OUT8_Mn9@258_g N_VSS_Mn9@258_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@259 N_OUT9_Mp9@259_d N_OUT8_Mp9@259_g N_VDD_Mp9@259_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@258 N_OUT9_Mp9@258_d N_OUT8_Mp9@258_g N_VDD_Mp9@258_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@257 N_OUT9_Mn9@257_d N_OUT8_Mn9@257_g N_VSS_Mn9@257_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@256 N_OUT9_Mn9@256_d N_OUT8_Mn9@256_g N_VSS_Mn9@256_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@257 N_OUT9_Mp9@257_d N_OUT8_Mp9@257_g N_VDD_Mp9@257_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@256 N_OUT9_Mp9@256_d N_OUT8_Mp9@256_g N_VDD_Mp9@256_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@255 N_OUT9_Mn9@255_d N_OUT8_Mn9@255_g N_VSS_Mn9@255_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@254 N_OUT9_Mn9@254_d N_OUT8_Mn9@254_g N_VSS_Mn9@254_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@255 N_OUT9_Mp9@255_d N_OUT8_Mp9@255_g N_VDD_Mp9@255_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@254 N_OUT9_Mp9@254_d N_OUT8_Mp9@254_g N_VDD_Mp9@254_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@253 N_OUT9_Mn9@253_d N_OUT8_Mn9@253_g N_VSS_Mn9@253_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@252 N_OUT9_Mn9@252_d N_OUT8_Mn9@252_g N_VSS_Mn9@252_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@253 N_OUT9_Mp9@253_d N_OUT8_Mp9@253_g N_VDD_Mp9@253_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@252 N_OUT9_Mp9@252_d N_OUT8_Mp9@252_g N_VDD_Mp9@252_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@251 N_OUT9_Mn9@251_d N_OUT8_Mn9@251_g N_VSS_Mn9@251_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@250 N_OUT9_Mn9@250_d N_OUT8_Mn9@250_g N_VSS_Mn9@250_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@251 N_OUT9_Mp9@251_d N_OUT8_Mp9@251_g N_VDD_Mp9@251_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@250 N_OUT9_Mp9@250_d N_OUT8_Mp9@250_g N_VDD_Mp9@250_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@249 N_OUT9_Mn9@249_d N_OUT8_Mn9@249_g N_VSS_Mn9@249_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@248 N_OUT9_Mn9@248_d N_OUT8_Mn9@248_g N_VSS_Mn9@248_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@249 N_OUT9_Mp9@249_d N_OUT8_Mp9@249_g N_VDD_Mp9@249_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@248 N_OUT9_Mp9@248_d N_OUT8_Mp9@248_g N_VDD_Mp9@248_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@247 N_OUT9_Mn9@247_d N_OUT8_Mn9@247_g N_VSS_Mn9@247_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@246 N_OUT9_Mn9@246_d N_OUT8_Mn9@246_g N_VSS_Mn9@246_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@247 N_OUT9_Mp9@247_d N_OUT8_Mp9@247_g N_VDD_Mp9@247_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@246 N_OUT9_Mp9@246_d N_OUT8_Mp9@246_g N_VDD_Mp9@246_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@245 N_OUT9_Mn9@245_d N_OUT8_Mn9@245_g N_VSS_Mn9@245_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@244 N_OUT9_Mn9@244_d N_OUT8_Mn9@244_g N_VSS_Mn9@244_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@245 N_OUT9_Mp9@245_d N_OUT8_Mp9@245_g N_VDD_Mp9@245_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@244 N_OUT9_Mp9@244_d N_OUT8_Mp9@244_g N_VDD_Mp9@244_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@243 N_OUT9_Mn9@243_d N_OUT8_Mn9@243_g N_VSS_Mn9@243_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@242 N_OUT9_Mn9@242_d N_OUT8_Mn9@242_g N_VSS_Mn9@242_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@243 N_OUT9_Mp9@243_d N_OUT8_Mp9@243_g N_VDD_Mp9@243_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@242 N_OUT9_Mp9@242_d N_OUT8_Mp9@242_g N_VDD_Mp9@242_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@241 N_OUT9_Mn9@241_d N_OUT8_Mn9@241_g N_VSS_Mn9@241_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@240 N_OUT9_Mn9@240_d N_OUT8_Mn9@240_g N_VSS_Mn9@240_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@241 N_OUT9_Mp9@241_d N_OUT8_Mp9@241_g N_VDD_Mp9@241_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@240 N_OUT9_Mp9@240_d N_OUT8_Mp9@240_g N_VDD_Mp9@240_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@239 N_OUT9_Mn9@239_d N_OUT8_Mn9@239_g N_VSS_Mn9@239_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@238 N_OUT9_Mn9@238_d N_OUT8_Mn9@238_g N_VSS_Mn9@238_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@239 N_OUT9_Mp9@239_d N_OUT8_Mp9@239_g N_VDD_Mp9@239_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@238 N_OUT9_Mp9@238_d N_OUT8_Mp9@238_g N_VDD_Mp9@238_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@237 N_OUT9_Mn9@237_d N_OUT8_Mn9@237_g N_VSS_Mn9@237_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@236 N_OUT9_Mn9@236_d N_OUT8_Mn9@236_g N_VSS_Mn9@236_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@237 N_OUT9_Mp9@237_d N_OUT8_Mp9@237_g N_VDD_Mp9@237_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@236 N_OUT9_Mp9@236_d N_OUT8_Mp9@236_g N_VDD_Mp9@236_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@235 N_OUT9_Mn9@235_d N_OUT8_Mn9@235_g N_VSS_Mn9@235_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@234 N_OUT9_Mn9@234_d N_OUT8_Mn9@234_g N_VSS_Mn9@234_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@235 N_OUT9_Mp9@235_d N_OUT8_Mp9@235_g N_VDD_Mp9@235_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@234 N_OUT9_Mp9@234_d N_OUT8_Mp9@234_g N_VDD_Mp9@234_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@233 N_OUT9_Mn9@233_d N_OUT8_Mn9@233_g N_VSS_Mn9@233_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@232 N_OUT9_Mn9@232_d N_OUT8_Mn9@232_g N_VSS_Mn9@232_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@233 N_OUT9_Mp9@233_d N_OUT8_Mp9@233_g N_VDD_Mp9@233_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@232 N_OUT9_Mp9@232_d N_OUT8_Mp9@232_g N_VDD_Mp9@232_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@231 N_OUT9_Mn9@231_d N_OUT8_Mn9@231_g N_VSS_Mn9@231_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@230 N_OUT9_Mn9@230_d N_OUT8_Mn9@230_g N_VSS_Mn9@230_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@231 N_OUT9_Mp9@231_d N_OUT8_Mp9@231_g N_VDD_Mp9@231_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@230 N_OUT9_Mp9@230_d N_OUT8_Mp9@230_g N_VDD_Mp9@230_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@229 N_OUT9_Mn9@229_d N_OUT8_Mn9@229_g N_VSS_Mn9@229_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@228 N_OUT9_Mn9@228_d N_OUT8_Mn9@228_g N_VSS_Mn9@228_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@229 N_OUT9_Mp9@229_d N_OUT8_Mp9@229_g N_VDD_Mp9@229_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@228 N_OUT9_Mp9@228_d N_OUT8_Mp9@228_g N_VDD_Mp9@228_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@227 N_OUT9_Mn9@227_d N_OUT8_Mn9@227_g N_VSS_Mn9@227_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@226 N_OUT9_Mn9@226_d N_OUT8_Mn9@226_g N_VSS_Mn9@226_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@227 N_OUT9_Mp9@227_d N_OUT8_Mp9@227_g N_VDD_Mp9@227_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@226 N_OUT9_Mp9@226_d N_OUT8_Mp9@226_g N_VDD_Mp9@226_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@225 N_OUT9_Mn9@225_d N_OUT8_Mn9@225_g N_VSS_Mn9@225_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@224 N_OUT9_Mn9@224_d N_OUT8_Mn9@224_g N_VSS_Mn9@224_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@225 N_OUT9_Mp9@225_d N_OUT8_Mp9@225_g N_VDD_Mp9@225_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@224 N_OUT9_Mp9@224_d N_OUT8_Mp9@224_g N_VDD_Mp9@224_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@223 N_OUT9_Mn9@223_d N_OUT8_Mn9@223_g N_VSS_Mn9@223_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@222 N_OUT9_Mn9@222_d N_OUT8_Mn9@222_g N_VSS_Mn9@222_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@223 N_OUT9_Mp9@223_d N_OUT8_Mp9@223_g N_VDD_Mp9@223_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@222 N_OUT9_Mp9@222_d N_OUT8_Mp9@222_g N_VDD_Mp9@222_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@221 N_OUT9_Mn9@221_d N_OUT8_Mn9@221_g N_VSS_Mn9@221_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@220 N_OUT9_Mn9@220_d N_OUT8_Mn9@220_g N_VSS_Mn9@220_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@221 N_OUT9_Mp9@221_d N_OUT8_Mp9@221_g N_VDD_Mp9@221_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@220 N_OUT9_Mp9@220_d N_OUT8_Mp9@220_g N_VDD_Mp9@220_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@219 N_OUT9_Mn9@219_d N_OUT8_Mn9@219_g N_VSS_Mn9@219_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@218 N_OUT9_Mn9@218_d N_OUT8_Mn9@218_g N_VSS_Mn9@218_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@219 N_OUT9_Mp9@219_d N_OUT8_Mp9@219_g N_VDD_Mp9@219_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@218 N_OUT9_Mp9@218_d N_OUT8_Mp9@218_g N_VDD_Mp9@218_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@217 N_OUT9_Mn9@217_d N_OUT8_Mn9@217_g N_VSS_Mn9@217_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@216 N_OUT9_Mn9@216_d N_OUT8_Mn9@216_g N_VSS_Mn9@216_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@217 N_OUT9_Mp9@217_d N_OUT8_Mp9@217_g N_VDD_Mp9@217_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@216 N_OUT9_Mp9@216_d N_OUT8_Mp9@216_g N_VDD_Mp9@216_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@215 N_OUT9_Mn9@215_d N_OUT8_Mn9@215_g N_VSS_Mn9@215_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@214 N_OUT9_Mn9@214_d N_OUT8_Mn9@214_g N_VSS_Mn9@214_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@215 N_OUT9_Mp9@215_d N_OUT8_Mp9@215_g N_VDD_Mp9@215_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@214 N_OUT9_Mp9@214_d N_OUT8_Mp9@214_g N_VDD_Mp9@214_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@213 N_OUT9_Mn9@213_d N_OUT8_Mn9@213_g N_VSS_Mn9@213_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@212 N_OUT9_Mn9@212_d N_OUT8_Mn9@212_g N_VSS_Mn9@212_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@213 N_OUT9_Mp9@213_d N_OUT8_Mp9@213_g N_VDD_Mp9@213_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@212 N_OUT9_Mp9@212_d N_OUT8_Mp9@212_g N_VDD_Mp9@212_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@211 N_OUT9_Mn9@211_d N_OUT8_Mn9@211_g N_VSS_Mn9@211_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@210 N_OUT9_Mn9@210_d N_OUT8_Mn9@210_g N_VSS_Mn9@210_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@211 N_OUT9_Mp9@211_d N_OUT8_Mp9@211_g N_VDD_Mp9@211_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@210 N_OUT9_Mp9@210_d N_OUT8_Mp9@210_g N_VDD_Mp9@210_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@209 N_OUT9_Mn9@209_d N_OUT8_Mn9@209_g N_VSS_Mn9@209_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@208 N_OUT9_Mn9@208_d N_OUT8_Mn9@208_g N_VSS_Mn9@208_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@209 N_OUT9_Mp9@209_d N_OUT8_Mp9@209_g N_VDD_Mp9@209_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@208 N_OUT9_Mp9@208_d N_OUT8_Mp9@208_g N_VDD_Mp9@208_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@207 N_OUT9_Mn9@207_d N_OUT8_Mn9@207_g N_VSS_Mn9@207_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@206 N_OUT9_Mn9@206_d N_OUT8_Mn9@206_g N_VSS_Mn9@206_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@207 N_OUT9_Mp9@207_d N_OUT8_Mp9@207_g N_VDD_Mp9@207_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@206 N_OUT9_Mp9@206_d N_OUT8_Mp9@206_g N_VDD_Mp9@206_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@205 N_OUT9_Mn9@205_d N_OUT8_Mn9@205_g N_VSS_Mn9@205_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@204 N_OUT9_Mn9@204_d N_OUT8_Mn9@204_g N_VSS_Mn9@204_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@205 N_OUT9_Mp9@205_d N_OUT8_Mp9@205_g N_VDD_Mp9@205_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@204 N_OUT9_Mp9@204_d N_OUT8_Mp9@204_g N_VDD_Mp9@204_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@203 N_OUT9_Mn9@203_d N_OUT8_Mn9@203_g N_VSS_Mn9@203_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@202 N_OUT9_Mn9@202_d N_OUT8_Mn9@202_g N_VSS_Mn9@202_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@203 N_OUT9_Mp9@203_d N_OUT8_Mp9@203_g N_VDD_Mp9@203_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@202 N_OUT9_Mp9@202_d N_OUT8_Mp9@202_g N_VDD_Mp9@202_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@201 N_OUT9_Mn9@201_d N_OUT8_Mn9@201_g N_VSS_Mn9@201_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@200 N_OUT9_Mn9@200_d N_OUT8_Mn9@200_g N_VSS_Mn9@200_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@201 N_OUT9_Mp9@201_d N_OUT8_Mp9@201_g N_VDD_Mp9@201_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@200 N_OUT9_Mp9@200_d N_OUT8_Mp9@200_g N_VDD_Mp9@200_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@199 N_OUT9_Mn9@199_d N_OUT8_Mn9@199_g N_VSS_Mn9@199_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@198 N_OUT9_Mn9@198_d N_OUT8_Mn9@198_g N_VSS_Mn9@198_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@199 N_OUT9_Mp9@199_d N_OUT8_Mp9@199_g N_VDD_Mp9@199_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@198 N_OUT9_Mp9@198_d N_OUT8_Mp9@198_g N_VDD_Mp9@198_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@197 N_OUT9_Mn9@197_d N_OUT8_Mn9@197_g N_VSS_Mn9@197_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@196 N_OUT9_Mn9@196_d N_OUT8_Mn9@196_g N_VSS_Mn9@196_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@197 N_OUT9_Mp9@197_d N_OUT8_Mp9@197_g N_VDD_Mp9@197_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@196 N_OUT9_Mp9@196_d N_OUT8_Mp9@196_g N_VDD_Mp9@196_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@195 N_OUT9_Mn9@195_d N_OUT8_Mn9@195_g N_VSS_Mn9@195_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@194 N_OUT9_Mn9@194_d N_OUT8_Mn9@194_g N_VSS_Mn9@194_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@195 N_OUT9_Mp9@195_d N_OUT8_Mp9@195_g N_VDD_Mp9@195_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@194 N_OUT9_Mp9@194_d N_OUT8_Mp9@194_g N_VDD_Mp9@194_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@193 N_OUT9_Mn9@193_d N_OUT8_Mn9@193_g N_VSS_Mn9@193_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@192 N_OUT9_Mn9@192_d N_OUT8_Mn9@192_g N_VSS_Mn9@192_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@193 N_OUT9_Mp9@193_d N_OUT8_Mp9@193_g N_VDD_Mp9@193_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@192 N_OUT9_Mp9@192_d N_OUT8_Mp9@192_g N_VDD_Mp9@192_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@191 N_OUT9_Mn9@191_d N_OUT8_Mn9@191_g N_VSS_Mn9@191_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@190 N_OUT9_Mn9@190_d N_OUT8_Mn9@190_g N_VSS_Mn9@190_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@191 N_OUT9_Mp9@191_d N_OUT8_Mp9@191_g N_VDD_Mp9@191_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@190 N_OUT9_Mp9@190_d N_OUT8_Mp9@190_g N_VDD_Mp9@190_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@189 N_OUT9_Mn9@189_d N_OUT8_Mn9@189_g N_VSS_Mn9@189_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@188 N_OUT9_Mn9@188_d N_OUT8_Mn9@188_g N_VSS_Mn9@188_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@189 N_OUT9_Mp9@189_d N_OUT8_Mp9@189_g N_VDD_Mp9@189_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@188 N_OUT9_Mp9@188_d N_OUT8_Mp9@188_g N_VDD_Mp9@188_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@187 N_OUT9_Mn9@187_d N_OUT8_Mn9@187_g N_VSS_Mn9@187_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@186 N_OUT9_Mn9@186_d N_OUT8_Mn9@186_g N_VSS_Mn9@186_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@187 N_OUT9_Mp9@187_d N_OUT8_Mp9@187_g N_VDD_Mp9@187_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@186 N_OUT9_Mp9@186_d N_OUT8_Mp9@186_g N_VDD_Mp9@186_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@185 N_OUT9_Mn9@185_d N_OUT8_Mn9@185_g N_VSS_Mn9@185_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@184 N_OUT9_Mn9@184_d N_OUT8_Mn9@184_g N_VSS_Mn9@184_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@185 N_OUT9_Mp9@185_d N_OUT8_Mp9@185_g N_VDD_Mp9@185_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@184 N_OUT9_Mp9@184_d N_OUT8_Mp9@184_g N_VDD_Mp9@184_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@183 N_OUT9_Mn9@183_d N_OUT8_Mn9@183_g N_VSS_Mn9@183_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@182 N_OUT9_Mn9@182_d N_OUT8_Mn9@182_g N_VSS_Mn9@182_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@183 N_OUT9_Mp9@183_d N_OUT8_Mp9@183_g N_VDD_Mp9@183_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@182 N_OUT9_Mp9@182_d N_OUT8_Mp9@182_g N_VDD_Mp9@182_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@181 N_OUT9_Mn9@181_d N_OUT8_Mn9@181_g N_VSS_Mn9@181_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@180 N_OUT9_Mn9@180_d N_OUT8_Mn9@180_g N_VSS_Mn9@180_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@181 N_OUT9_Mp9@181_d N_OUT8_Mp9@181_g N_VDD_Mp9@181_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@180 N_OUT9_Mp9@180_d N_OUT8_Mp9@180_g N_VDD_Mp9@180_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@179 N_OUT9_Mn9@179_d N_OUT8_Mn9@179_g N_VSS_Mn9@179_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@178 N_OUT9_Mn9@178_d N_OUT8_Mn9@178_g N_VSS_Mn9@178_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@179 N_OUT9_Mp9@179_d N_OUT8_Mp9@179_g N_VDD_Mp9@179_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@178 N_OUT9_Mp9@178_d N_OUT8_Mp9@178_g N_VDD_Mp9@178_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@177 N_OUT9_Mn9@177_d N_OUT8_Mn9@177_g N_VSS_Mn9@177_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@176 N_OUT9_Mn9@176_d N_OUT8_Mn9@176_g N_VSS_Mn9@176_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@177 N_OUT9_Mp9@177_d N_OUT8_Mp9@177_g N_VDD_Mp9@177_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@176 N_OUT9_Mp9@176_d N_OUT8_Mp9@176_g N_VDD_Mp9@176_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@175 N_OUT9_Mn9@175_d N_OUT8_Mn9@175_g N_VSS_Mn9@175_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@174 N_OUT9_Mn9@174_d N_OUT8_Mn9@174_g N_VSS_Mn9@174_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@175 N_OUT9_Mp9@175_d N_OUT8_Mp9@175_g N_VDD_Mp9@175_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@174 N_OUT9_Mp9@174_d N_OUT8_Mp9@174_g N_VDD_Mp9@174_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@173 N_OUT9_Mn9@173_d N_OUT8_Mn9@173_g N_VSS_Mn9@173_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@172 N_OUT9_Mn9@172_d N_OUT8_Mn9@172_g N_VSS_Mn9@172_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@173 N_OUT9_Mp9@173_d N_OUT8_Mp9@173_g N_VDD_Mp9@173_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@172 N_OUT9_Mp9@172_d N_OUT8_Mp9@172_g N_VDD_Mp9@172_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@171 N_OUT9_Mn9@171_d N_OUT8_Mn9@171_g N_VSS_Mn9@171_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@170 N_OUT9_Mn9@170_d N_OUT8_Mn9@170_g N_VSS_Mn9@170_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@171 N_OUT9_Mp9@171_d N_OUT8_Mp9@171_g N_VDD_Mp9@171_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@170 N_OUT9_Mp9@170_d N_OUT8_Mp9@170_g N_VDD_Mp9@170_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@169 N_OUT9_Mn9@169_d N_OUT8_Mn9@169_g N_VSS_Mn9@169_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@168 N_OUT9_Mn9@168_d N_OUT8_Mn9@168_g N_VSS_Mn9@168_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@169 N_OUT9_Mp9@169_d N_OUT8_Mp9@169_g N_VDD_Mp9@169_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@168 N_OUT9_Mp9@168_d N_OUT8_Mp9@168_g N_VDD_Mp9@168_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@167 N_OUT9_Mn9@167_d N_OUT8_Mn9@167_g N_VSS_Mn9@167_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@166 N_OUT9_Mn9@166_d N_OUT8_Mn9@166_g N_VSS_Mn9@166_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@167 N_OUT9_Mp9@167_d N_OUT8_Mp9@167_g N_VDD_Mp9@167_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@166 N_OUT9_Mp9@166_d N_OUT8_Mp9@166_g N_VDD_Mp9@166_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@165 N_OUT9_Mn9@165_d N_OUT8_Mn9@165_g N_VSS_Mn9@165_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@164 N_OUT9_Mn9@164_d N_OUT8_Mn9@164_g N_VSS_Mn9@164_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@165 N_OUT9_Mp9@165_d N_OUT8_Mp9@165_g N_VDD_Mp9@165_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@164 N_OUT9_Mp9@164_d N_OUT8_Mp9@164_g N_VDD_Mp9@164_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@163 N_OUT9_Mn9@163_d N_OUT8_Mn9@163_g N_VSS_Mn9@163_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@162 N_OUT9_Mn9@162_d N_OUT8_Mn9@162_g N_VSS_Mn9@162_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@163 N_OUT9_Mp9@163_d N_OUT8_Mp9@163_g N_VDD_Mp9@163_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@162 N_OUT9_Mp9@162_d N_OUT8_Mp9@162_g N_VDD_Mp9@162_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@161 N_OUT9_Mn9@161_d N_OUT8_Mn9@161_g N_VSS_Mn9@161_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@160 N_OUT9_Mn9@160_d N_OUT8_Mn9@160_g N_VSS_Mn9@160_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@161 N_OUT9_Mp9@161_d N_OUT8_Mp9@161_g N_VDD_Mp9@161_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@160 N_OUT9_Mp9@160_d N_OUT8_Mp9@160_g N_VDD_Mp9@160_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@159 N_OUT9_Mn9@159_d N_OUT8_Mn9@159_g N_VSS_Mn9@159_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@158 N_OUT9_Mn9@158_d N_OUT8_Mn9@158_g N_VSS_Mn9@158_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@159 N_OUT9_Mp9@159_d N_OUT8_Mp9@159_g N_VDD_Mp9@159_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@158 N_OUT9_Mp9@158_d N_OUT8_Mp9@158_g N_VDD_Mp9@158_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@157 N_OUT9_Mn9@157_d N_OUT8_Mn9@157_g N_VSS_Mn9@157_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@156 N_OUT9_Mn9@156_d N_OUT8_Mn9@156_g N_VSS_Mn9@156_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@157 N_OUT9_Mp9@157_d N_OUT8_Mp9@157_g N_VDD_Mp9@157_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@156 N_OUT9_Mp9@156_d N_OUT8_Mp9@156_g N_VDD_Mp9@156_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@155 N_OUT9_Mn9@155_d N_OUT8_Mn9@155_g N_VSS_Mn9@155_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@154 N_OUT9_Mn9@154_d N_OUT8_Mn9@154_g N_VSS_Mn9@154_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@155 N_OUT9_Mp9@155_d N_OUT8_Mp9@155_g N_VDD_Mp9@155_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@154 N_OUT9_Mp9@154_d N_OUT8_Mp9@154_g N_VDD_Mp9@154_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@153 N_OUT9_Mn9@153_d N_OUT8_Mn9@153_g N_VSS_Mn9@153_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@152 N_OUT9_Mn9@152_d N_OUT8_Mn9@152_g N_VSS_Mn9@152_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@153 N_OUT9_Mp9@153_d N_OUT8_Mp9@153_g N_VDD_Mp9@153_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@152 N_OUT9_Mp9@152_d N_OUT8_Mp9@152_g N_VDD_Mp9@152_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@151 N_OUT9_Mn9@151_d N_OUT8_Mn9@151_g N_VSS_Mn9@151_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@150 N_OUT9_Mn9@150_d N_OUT8_Mn9@150_g N_VSS_Mn9@150_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@151 N_OUT9_Mp9@151_d N_OUT8_Mp9@151_g N_VDD_Mp9@151_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@150 N_OUT9_Mp9@150_d N_OUT8_Mp9@150_g N_VDD_Mp9@150_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@149 N_OUT9_Mn9@149_d N_OUT8_Mn9@149_g N_VSS_Mn9@149_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@148 N_OUT9_Mn9@148_d N_OUT8_Mn9@148_g N_VSS_Mn9@148_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@149 N_OUT9_Mp9@149_d N_OUT8_Mp9@149_g N_VDD_Mp9@149_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@148 N_OUT9_Mp9@148_d N_OUT8_Mp9@148_g N_VDD_Mp9@148_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@147 N_OUT9_Mn9@147_d N_OUT8_Mn9@147_g N_VSS_Mn9@147_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@146 N_OUT9_Mn9@146_d N_OUT8_Mn9@146_g N_VSS_Mn9@146_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@147 N_OUT9_Mp9@147_d N_OUT8_Mp9@147_g N_VDD_Mp9@147_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@146 N_OUT9_Mp9@146_d N_OUT8_Mp9@146_g N_VDD_Mp9@146_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@145 N_OUT9_Mn9@145_d N_OUT8_Mn9@145_g N_VSS_Mn9@145_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@144 N_OUT9_Mn9@144_d N_OUT8_Mn9@144_g N_VSS_Mn9@144_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@145 N_OUT9_Mp9@145_d N_OUT8_Mp9@145_g N_VDD_Mp9@145_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@144 N_OUT9_Mp9@144_d N_OUT8_Mp9@144_g N_VDD_Mp9@144_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@143 N_OUT9_Mn9@143_d N_OUT8_Mn9@143_g N_VSS_Mn9@143_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@142 N_OUT9_Mn9@142_d N_OUT8_Mn9@142_g N_VSS_Mn9@142_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@143 N_OUT9_Mp9@143_d N_OUT8_Mp9@143_g N_VDD_Mp9@143_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@142 N_OUT9_Mp9@142_d N_OUT8_Mp9@142_g N_VDD_Mp9@142_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@141 N_OUT9_Mn9@141_d N_OUT8_Mn9@141_g N_VSS_Mn9@141_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@140 N_OUT9_Mn9@140_d N_OUT8_Mn9@140_g N_VSS_Mn9@140_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@141 N_OUT9_Mp9@141_d N_OUT8_Mp9@141_g N_VDD_Mp9@141_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@140 N_OUT9_Mp9@140_d N_OUT8_Mp9@140_g N_VDD_Mp9@140_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@139 N_OUT9_Mn9@139_d N_OUT8_Mn9@139_g N_VSS_Mn9@139_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@138 N_OUT9_Mn9@138_d N_OUT8_Mn9@138_g N_VSS_Mn9@138_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@139 N_OUT9_Mp9@139_d N_OUT8_Mp9@139_g N_VDD_Mp9@139_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@138 N_OUT9_Mp9@138_d N_OUT8_Mp9@138_g N_VDD_Mp9@138_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@137 N_OUT9_Mn9@137_d N_OUT8_Mn9@137_g N_VSS_Mn9@137_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@136 N_OUT9_Mn9@136_d N_OUT8_Mn9@136_g N_VSS_Mn9@136_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@137 N_OUT9_Mp9@137_d N_OUT8_Mp9@137_g N_VDD_Mp9@137_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@136 N_OUT9_Mp9@136_d N_OUT8_Mp9@136_g N_VDD_Mp9@136_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@135 N_OUT9_Mn9@135_d N_OUT8_Mn9@135_g N_VSS_Mn9@135_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@134 N_OUT9_Mn9@134_d N_OUT8_Mn9@134_g N_VSS_Mn9@134_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@135 N_OUT9_Mp9@135_d N_OUT8_Mp9@135_g N_VDD_Mp9@135_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@134 N_OUT9_Mp9@134_d N_OUT8_Mp9@134_g N_VDD_Mp9@134_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@133 N_OUT9_Mn9@133_d N_OUT8_Mn9@133_g N_VSS_Mn9@133_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@132 N_OUT9_Mn9@132_d N_OUT8_Mn9@132_g N_VSS_Mn9@132_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@133 N_OUT9_Mp9@133_d N_OUT8_Mp9@133_g N_VDD_Mp9@133_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@132 N_OUT9_Mp9@132_d N_OUT8_Mp9@132_g N_VDD_Mp9@132_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@131 N_OUT9_Mn9@131_d N_OUT8_Mn9@131_g N_VSS_Mn9@131_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@130 N_OUT9_Mn9@130_d N_OUT8_Mn9@130_g N_VSS_Mn9@130_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@131 N_OUT9_Mp9@131_d N_OUT8_Mp9@131_g N_VDD_Mp9@131_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@130 N_OUT9_Mp9@130_d N_OUT8_Mp9@130_g N_VDD_Mp9@130_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@129 N_OUT9_Mn9@129_d N_OUT8_Mn9@129_g N_VSS_Mn9@129_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@128 N_OUT9_Mn9@128_d N_OUT8_Mn9@128_g N_VSS_Mn9@128_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@129 N_OUT9_Mp9@129_d N_OUT8_Mp9@129_g N_VDD_Mp9@129_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@128 N_OUT9_Mp9@128_d N_OUT8_Mp9@128_g N_VDD_Mp9@128_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@127 N_OUT9_Mn9@127_d N_OUT8_Mn9@127_g N_VSS_Mn9@127_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@126 N_OUT9_Mn9@126_d N_OUT8_Mn9@126_g N_VSS_Mn9@126_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@127 N_OUT9_Mp9@127_d N_OUT8_Mp9@127_g N_VDD_Mp9@127_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@126 N_OUT9_Mp9@126_d N_OUT8_Mp9@126_g N_VDD_Mp9@126_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@125 N_OUT9_Mn9@125_d N_OUT8_Mn9@125_g N_VSS_Mn9@125_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@124 N_OUT9_Mn9@124_d N_OUT8_Mn9@124_g N_VSS_Mn9@124_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@125 N_OUT9_Mp9@125_d N_OUT8_Mp9@125_g N_VDD_Mp9@125_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@124 N_OUT9_Mp9@124_d N_OUT8_Mp9@124_g N_VDD_Mp9@124_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@123 N_OUT9_Mn9@123_d N_OUT8_Mn9@123_g N_VSS_Mn9@123_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@122 N_OUT9_Mn9@122_d N_OUT8_Mn9@122_g N_VSS_Mn9@122_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@123 N_OUT9_Mp9@123_d N_OUT8_Mp9@123_g N_VDD_Mp9@123_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@122 N_OUT9_Mp9@122_d N_OUT8_Mp9@122_g N_VDD_Mp9@122_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@121 N_OUT9_Mn9@121_d N_OUT8_Mn9@121_g N_VSS_Mn9@121_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@120 N_OUT9_Mn9@120_d N_OUT8_Mn9@120_g N_VSS_Mn9@120_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@121 N_OUT9_Mp9@121_d N_OUT8_Mp9@121_g N_VDD_Mp9@121_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@120 N_OUT9_Mp9@120_d N_OUT8_Mp9@120_g N_VDD_Mp9@120_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@119 N_OUT9_Mn9@119_d N_OUT8_Mn9@119_g N_VSS_Mn9@119_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@118 N_OUT9_Mn9@118_d N_OUT8_Mn9@118_g N_VSS_Mn9@118_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@119 N_OUT9_Mp9@119_d N_OUT8_Mp9@119_g N_VDD_Mp9@119_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@118 N_OUT9_Mp9@118_d N_OUT8_Mp9@118_g N_VDD_Mp9@118_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@117 N_OUT9_Mn9@117_d N_OUT8_Mn9@117_g N_VSS_Mn9@117_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@116 N_OUT9_Mn9@116_d N_OUT8_Mn9@116_g N_VSS_Mn9@116_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@117 N_OUT9_Mp9@117_d N_OUT8_Mp9@117_g N_VDD_Mp9@117_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@116 N_OUT9_Mp9@116_d N_OUT8_Mp9@116_g N_VDD_Mp9@116_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@115 N_OUT9_Mn9@115_d N_OUT8_Mn9@115_g N_VSS_Mn9@115_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@114 N_OUT9_Mn9@114_d N_OUT8_Mn9@114_g N_VSS_Mn9@114_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@115 N_OUT9_Mp9@115_d N_OUT8_Mp9@115_g N_VDD_Mp9@115_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@114 N_OUT9_Mp9@114_d N_OUT8_Mp9@114_g N_VDD_Mp9@114_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@113 N_OUT9_Mn9@113_d N_OUT8_Mn9@113_g N_VSS_Mn9@113_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@112 N_OUT9_Mn9@112_d N_OUT8_Mn9@112_g N_VSS_Mn9@112_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@113 N_OUT9_Mp9@113_d N_OUT8_Mp9@113_g N_VDD_Mp9@113_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@112 N_OUT9_Mp9@112_d N_OUT8_Mp9@112_g N_VDD_Mp9@112_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@111 N_OUT9_Mn9@111_d N_OUT8_Mn9@111_g N_VSS_Mn9@111_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@110 N_OUT9_Mn9@110_d N_OUT8_Mn9@110_g N_VSS_Mn9@110_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@111 N_OUT9_Mp9@111_d N_OUT8_Mp9@111_g N_VDD_Mp9@111_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@110 N_OUT9_Mp9@110_d N_OUT8_Mp9@110_g N_VDD_Mp9@110_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@109 N_OUT9_Mn9@109_d N_OUT8_Mn9@109_g N_VSS_Mn9@109_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@108 N_OUT9_Mn9@108_d N_OUT8_Mn9@108_g N_VSS_Mn9@108_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@109 N_OUT9_Mp9@109_d N_OUT8_Mp9@109_g N_VDD_Mp9@109_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@108 N_OUT9_Mp9@108_d N_OUT8_Mp9@108_g N_VDD_Mp9@108_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@107 N_OUT9_Mn9@107_d N_OUT8_Mn9@107_g N_VSS_Mn9@107_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@106 N_OUT9_Mn9@106_d N_OUT8_Mn9@106_g N_VSS_Mn9@106_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@107 N_OUT9_Mp9@107_d N_OUT8_Mp9@107_g N_VDD_Mp9@107_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@106 N_OUT9_Mp9@106_d N_OUT8_Mp9@106_g N_VDD_Mp9@106_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@105 N_OUT9_Mn9@105_d N_OUT8_Mn9@105_g N_VSS_Mn9@105_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@104 N_OUT9_Mn9@104_d N_OUT8_Mn9@104_g N_VSS_Mn9@104_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@105 N_OUT9_Mp9@105_d N_OUT8_Mp9@105_g N_VDD_Mp9@105_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@104 N_OUT9_Mp9@104_d N_OUT8_Mp9@104_g N_VDD_Mp9@104_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@103 N_OUT9_Mn9@103_d N_OUT8_Mn9@103_g N_VSS_Mn9@103_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@102 N_OUT9_Mn9@102_d N_OUT8_Mn9@102_g N_VSS_Mn9@102_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@103 N_OUT9_Mp9@103_d N_OUT8_Mp9@103_g N_VDD_Mp9@103_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@102 N_OUT9_Mp9@102_d N_OUT8_Mp9@102_g N_VDD_Mp9@102_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@101 N_OUT9_Mn9@101_d N_OUT8_Mn9@101_g N_VSS_Mn9@101_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@100 N_OUT9_Mn9@100_d N_OUT8_Mn9@100_g N_VSS_Mn9@100_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@101 N_OUT9_Mp9@101_d N_OUT8_Mp9@101_g N_VDD_Mp9@101_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@100 N_OUT9_Mp9@100_d N_OUT8_Mp9@100_g N_VDD_Mp9@100_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@99 N_OUT9_Mn9@99_d N_OUT8_Mn9@99_g N_VSS_Mn9@99_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@98 N_OUT9_Mn9@98_d N_OUT8_Mn9@98_g N_VSS_Mn9@98_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@99 N_OUT9_Mp9@99_d N_OUT8_Mp9@99_g N_VDD_Mp9@99_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@98 N_OUT9_Mp9@98_d N_OUT8_Mp9@98_g N_VDD_Mp9@98_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@97 N_OUT9_Mn9@97_d N_OUT8_Mn9@97_g N_VSS_Mn9@97_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@96 N_OUT9_Mn9@96_d N_OUT8_Mn9@96_g N_VSS_Mn9@96_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@97 N_OUT9_Mp9@97_d N_OUT8_Mp9@97_g N_VDD_Mp9@97_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@96 N_OUT9_Mp9@96_d N_OUT8_Mp9@96_g N_VDD_Mp9@96_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@95 N_OUT9_Mn9@95_d N_OUT8_Mn9@95_g N_VSS_Mn9@95_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@94 N_OUT9_Mn9@94_d N_OUT8_Mn9@94_g N_VSS_Mn9@94_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@95 N_OUT9_Mp9@95_d N_OUT8_Mp9@95_g N_VDD_Mp9@95_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@94 N_OUT9_Mp9@94_d N_OUT8_Mp9@94_g N_VDD_Mp9@94_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@93 N_OUT9_Mn9@93_d N_OUT8_Mn9@93_g N_VSS_Mn9@93_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@92 N_OUT9_Mn9@92_d N_OUT8_Mn9@92_g N_VSS_Mn9@92_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@93 N_OUT9_Mp9@93_d N_OUT8_Mp9@93_g N_VDD_Mp9@93_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@92 N_OUT9_Mp9@92_d N_OUT8_Mp9@92_g N_VDD_Mp9@92_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@91 N_OUT9_Mn9@91_d N_OUT8_Mn9@91_g N_VSS_Mn9@91_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@90 N_OUT9_Mn9@90_d N_OUT8_Mn9@90_g N_VSS_Mn9@90_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@91 N_OUT9_Mp9@91_d N_OUT8_Mp9@91_g N_VDD_Mp9@91_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@90 N_OUT9_Mp9@90_d N_OUT8_Mp9@90_g N_VDD_Mp9@90_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@89 N_OUT9_Mn9@89_d N_OUT8_Mn9@89_g N_VSS_Mn9@89_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@88 N_OUT9_Mn9@88_d N_OUT8_Mn9@88_g N_VSS_Mn9@88_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@89 N_OUT9_Mp9@89_d N_OUT8_Mp9@89_g N_VDD_Mp9@89_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@88 N_OUT9_Mp9@88_d N_OUT8_Mp9@88_g N_VDD_Mp9@88_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@87 N_OUT9_Mn9@87_d N_OUT8_Mn9@87_g N_VSS_Mn9@87_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@86 N_OUT9_Mn9@86_d N_OUT8_Mn9@86_g N_VSS_Mn9@86_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@87 N_OUT9_Mp9@87_d N_OUT8_Mp9@87_g N_VDD_Mp9@87_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@86 N_OUT9_Mp9@86_d N_OUT8_Mp9@86_g N_VDD_Mp9@86_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@85 N_OUT9_Mn9@85_d N_OUT8_Mn9@85_g N_VSS_Mn9@85_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@84 N_OUT9_Mn9@84_d N_OUT8_Mn9@84_g N_VSS_Mn9@84_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@85 N_OUT9_Mp9@85_d N_OUT8_Mp9@85_g N_VDD_Mp9@85_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@84 N_OUT9_Mp9@84_d N_OUT8_Mp9@84_g N_VDD_Mp9@84_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@83 N_OUT9_Mn9@83_d N_OUT8_Mn9@83_g N_VSS_Mn9@83_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@82 N_OUT9_Mn9@82_d N_OUT8_Mn9@82_g N_VSS_Mn9@82_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@83 N_OUT9_Mp9@83_d N_OUT8_Mp9@83_g N_VDD_Mp9@83_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@82 N_OUT9_Mp9@82_d N_OUT8_Mp9@82_g N_VDD_Mp9@82_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@81 N_OUT9_Mn9@81_d N_OUT8_Mn9@81_g N_VSS_Mn9@81_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@80 N_OUT9_Mn9@80_d N_OUT8_Mn9@80_g N_VSS_Mn9@80_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@81 N_OUT9_Mp9@81_d N_OUT8_Mp9@81_g N_VDD_Mp9@81_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@80 N_OUT9_Mp9@80_d N_OUT8_Mp9@80_g N_VDD_Mp9@80_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@79 N_OUT9_Mn9@79_d N_OUT8_Mn9@79_g N_VSS_Mn9@79_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@78 N_OUT9_Mn9@78_d N_OUT8_Mn9@78_g N_VSS_Mn9@78_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@79 N_OUT9_Mp9@79_d N_OUT8_Mp9@79_g N_VDD_Mp9@79_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@78 N_OUT9_Mp9@78_d N_OUT8_Mp9@78_g N_VDD_Mp9@78_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@77 N_OUT9_Mn9@77_d N_OUT8_Mn9@77_g N_VSS_Mn9@77_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@76 N_OUT9_Mn9@76_d N_OUT8_Mn9@76_g N_VSS_Mn9@76_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@77 N_OUT9_Mp9@77_d N_OUT8_Mp9@77_g N_VDD_Mp9@77_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@76 N_OUT9_Mp9@76_d N_OUT8_Mp9@76_g N_VDD_Mp9@76_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@75 N_OUT9_Mn9@75_d N_OUT8_Mn9@75_g N_VSS_Mn9@75_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@74 N_OUT9_Mn9@74_d N_OUT8_Mn9@74_g N_VSS_Mn9@74_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@75 N_OUT9_Mp9@75_d N_OUT8_Mp9@75_g N_VDD_Mp9@75_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@74 N_OUT9_Mp9@74_d N_OUT8_Mp9@74_g N_VDD_Mp9@74_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@73 N_OUT9_Mn9@73_d N_OUT8_Mn9@73_g N_VSS_Mn9@73_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@72 N_OUT9_Mn9@72_d N_OUT8_Mn9@72_g N_VSS_Mn9@72_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@73 N_OUT9_Mp9@73_d N_OUT8_Mp9@73_g N_VDD_Mp9@73_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@72 N_OUT9_Mp9@72_d N_OUT8_Mp9@72_g N_VDD_Mp9@72_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@71 N_OUT9_Mn9@71_d N_OUT8_Mn9@71_g N_VSS_Mn9@71_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@70 N_OUT9_Mn9@70_d N_OUT8_Mn9@70_g N_VSS_Mn9@70_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@71 N_OUT9_Mp9@71_d N_OUT8_Mp9@71_g N_VDD_Mp9@71_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@70 N_OUT9_Mp9@70_d N_OUT8_Mp9@70_g N_VDD_Mp9@70_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@69 N_OUT9_Mn9@69_d N_OUT8_Mn9@69_g N_VSS_Mn9@69_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@68 N_OUT9_Mn9@68_d N_OUT8_Mn9@68_g N_VSS_Mn9@68_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@69 N_OUT9_Mp9@69_d N_OUT8_Mp9@69_g N_VDD_Mp9@69_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@68 N_OUT9_Mp9@68_d N_OUT8_Mp9@68_g N_VDD_Mp9@68_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@67 N_OUT9_Mn9@67_d N_OUT8_Mn9@67_g N_VSS_Mn9@67_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@66 N_OUT9_Mn9@66_d N_OUT8_Mn9@66_g N_VSS_Mn9@66_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@67 N_OUT9_Mp9@67_d N_OUT8_Mp9@67_g N_VDD_Mp9@67_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@66 N_OUT9_Mp9@66_d N_OUT8_Mp9@66_g N_VDD_Mp9@66_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@65 N_OUT9_Mn9@65_d N_OUT8_Mn9@65_g N_VSS_Mn9@65_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@64 N_OUT9_Mn9@64_d N_OUT8_Mn9@64_g N_VSS_Mn9@64_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@65 N_OUT9_Mp9@65_d N_OUT8_Mp9@65_g N_VDD_Mp9@65_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@64 N_OUT9_Mp9@64_d N_OUT8_Mp9@64_g N_VDD_Mp9@64_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@63 N_OUT9_Mn9@63_d N_OUT8_Mn9@63_g N_VSS_Mn9@63_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@62 N_OUT9_Mn9@62_d N_OUT8_Mn9@62_g N_VSS_Mn9@62_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@63 N_OUT9_Mp9@63_d N_OUT8_Mp9@63_g N_VDD_Mp9@63_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@62 N_OUT9_Mp9@62_d N_OUT8_Mp9@62_g N_VDD_Mp9@62_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@61 N_OUT9_Mn9@61_d N_OUT8_Mn9@61_g N_VSS_Mn9@61_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@60 N_OUT9_Mn9@60_d N_OUT8_Mn9@60_g N_VSS_Mn9@60_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@61 N_OUT9_Mp9@61_d N_OUT8_Mp9@61_g N_VDD_Mp9@61_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@60 N_OUT9_Mp9@60_d N_OUT8_Mp9@60_g N_VDD_Mp9@60_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@59 N_OUT9_Mn9@59_d N_OUT8_Mn9@59_g N_VSS_Mn9@59_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@58 N_OUT9_Mn9@58_d N_OUT8_Mn9@58_g N_VSS_Mn9@58_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@59 N_OUT9_Mp9@59_d N_OUT8_Mp9@59_g N_VDD_Mp9@59_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@58 N_OUT9_Mp9@58_d N_OUT8_Mp9@58_g N_VDD_Mp9@58_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@57 N_OUT9_Mn9@57_d N_OUT8_Mn9@57_g N_VSS_Mn9@57_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@56 N_OUT9_Mn9@56_d N_OUT8_Mn9@56_g N_VSS_Mn9@56_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@57 N_OUT9_Mp9@57_d N_OUT8_Mp9@57_g N_VDD_Mp9@57_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@56 N_OUT9_Mp9@56_d N_OUT8_Mp9@56_g N_VDD_Mp9@56_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@55 N_OUT9_Mn9@55_d N_OUT8_Mn9@55_g N_VSS_Mn9@55_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@54 N_OUT9_Mn9@54_d N_OUT8_Mn9@54_g N_VSS_Mn9@54_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@55 N_OUT9_Mp9@55_d N_OUT8_Mp9@55_g N_VDD_Mp9@55_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@54 N_OUT9_Mp9@54_d N_OUT8_Mp9@54_g N_VDD_Mp9@54_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@53 N_OUT9_Mn9@53_d N_OUT8_Mn9@53_g N_VSS_Mn9@53_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@52 N_OUT9_Mn9@52_d N_OUT8_Mn9@52_g N_VSS_Mn9@52_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@53 N_OUT9_Mp9@53_d N_OUT8_Mp9@53_g N_VDD_Mp9@53_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@52 N_OUT9_Mp9@52_d N_OUT8_Mp9@52_g N_VDD_Mp9@52_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@51 N_OUT9_Mn9@51_d N_OUT8_Mn9@51_g N_VSS_Mn9@51_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@50 N_OUT9_Mn9@50_d N_OUT8_Mn9@50_g N_VSS_Mn9@50_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@51 N_OUT9_Mp9@51_d N_OUT8_Mp9@51_g N_VDD_Mp9@51_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@50 N_OUT9_Mp9@50_d N_OUT8_Mp9@50_g N_VDD_Mp9@50_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@49 N_OUT9_Mn9@49_d N_OUT8_Mn9@49_g N_VSS_Mn9@49_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@48 N_OUT9_Mn9@48_d N_OUT8_Mn9@48_g N_VSS_Mn9@48_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@49 N_OUT9_Mp9@49_d N_OUT8_Mp9@49_g N_VDD_Mp9@49_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@48 N_OUT9_Mp9@48_d N_OUT8_Mp9@48_g N_VDD_Mp9@48_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@47 N_OUT9_Mn9@47_d N_OUT8_Mn9@47_g N_VSS_Mn9@47_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@46 N_OUT9_Mn9@46_d N_OUT8_Mn9@46_g N_VSS_Mn9@46_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@47 N_OUT9_Mp9@47_d N_OUT8_Mp9@47_g N_VDD_Mp9@47_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@46 N_OUT9_Mp9@46_d N_OUT8_Mp9@46_g N_VDD_Mp9@46_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@45 N_OUT9_Mn9@45_d N_OUT8_Mn9@45_g N_VSS_Mn9@45_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@44 N_OUT9_Mn9@44_d N_OUT8_Mn9@44_g N_VSS_Mn9@44_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@45 N_OUT9_Mp9@45_d N_OUT8_Mp9@45_g N_VDD_Mp9@45_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@44 N_OUT9_Mp9@44_d N_OUT8_Mp9@44_g N_VDD_Mp9@44_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@43 N_OUT9_Mn9@43_d N_OUT8_Mn9@43_g N_VSS_Mn9@43_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@42 N_OUT9_Mn9@42_d N_OUT8_Mn9@42_g N_VSS_Mn9@42_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@43 N_OUT9_Mp9@43_d N_OUT8_Mp9@43_g N_VDD_Mp9@43_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@42 N_OUT9_Mp9@42_d N_OUT8_Mp9@42_g N_VDD_Mp9@42_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@41 N_OUT9_Mn9@41_d N_OUT8_Mn9@41_g N_VSS_Mn9@41_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@40 N_OUT9_Mn9@40_d N_OUT8_Mn9@40_g N_VSS_Mn9@40_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@41 N_OUT9_Mp9@41_d N_OUT8_Mp9@41_g N_VDD_Mp9@41_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@40 N_OUT9_Mp9@40_d N_OUT8_Mp9@40_g N_VDD_Mp9@40_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@39 N_OUT9_Mn9@39_d N_OUT8_Mn9@39_g N_VSS_Mn9@39_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@38 N_OUT9_Mn9@38_d N_OUT8_Mn9@38_g N_VSS_Mn9@38_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@39 N_OUT9_Mp9@39_d N_OUT8_Mp9@39_g N_VDD_Mp9@39_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@38 N_OUT9_Mp9@38_d N_OUT8_Mp9@38_g N_VDD_Mp9@38_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@37 N_OUT9_Mn9@37_d N_OUT8_Mn9@37_g N_VSS_Mn9@37_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@36 N_OUT9_Mn9@36_d N_OUT8_Mn9@36_g N_VSS_Mn9@36_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@37 N_OUT9_Mp9@37_d N_OUT8_Mp9@37_g N_VDD_Mp9@37_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@36 N_OUT9_Mp9@36_d N_OUT8_Mp9@36_g N_VDD_Mp9@36_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@35 N_OUT9_Mn9@35_d N_OUT8_Mn9@35_g N_VSS_Mn9@35_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@34 N_OUT9_Mn9@34_d N_OUT8_Mn9@34_g N_VSS_Mn9@34_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@35 N_OUT9_Mp9@35_d N_OUT8_Mp9@35_g N_VDD_Mp9@35_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@34 N_OUT9_Mp9@34_d N_OUT8_Mp9@34_g N_VDD_Mp9@34_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@33 N_OUT9_Mn9@33_d N_OUT8_Mn9@33_g N_VSS_Mn9@33_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@32 N_OUT9_Mn9@32_d N_OUT8_Mn9@32_g N_VSS_Mn9@32_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@33 N_OUT9_Mp9@33_d N_OUT8_Mp9@33_g N_VDD_Mp9@33_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@32 N_OUT9_Mp9@32_d N_OUT8_Mp9@32_g N_VDD_Mp9@32_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@31 N_OUT9_Mn9@31_d N_OUT8_Mn9@31_g N_VSS_Mn9@31_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@30 N_OUT9_Mn9@30_d N_OUT8_Mn9@30_g N_VSS_Mn9@30_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@31 N_OUT9_Mp9@31_d N_OUT8_Mp9@31_g N_VDD_Mp9@31_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@30 N_OUT9_Mp9@30_d N_OUT8_Mp9@30_g N_VDD_Mp9@30_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@29 N_OUT9_Mn9@29_d N_OUT8_Mn9@29_g N_VSS_Mn9@29_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@28 N_OUT9_Mn9@28_d N_OUT8_Mn9@28_g N_VSS_Mn9@28_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@29 N_OUT9_Mp9@29_d N_OUT8_Mp9@29_g N_VDD_Mp9@29_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@28 N_OUT9_Mp9@28_d N_OUT8_Mp9@28_g N_VDD_Mp9@28_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@27 N_OUT9_Mn9@27_d N_OUT8_Mn9@27_g N_VSS_Mn9@27_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@26 N_OUT9_Mn9@26_d N_OUT8_Mn9@26_g N_VSS_Mn9@26_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@27 N_OUT9_Mp9@27_d N_OUT8_Mp9@27_g N_VDD_Mp9@27_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@26 N_OUT9_Mp9@26_d N_OUT8_Mp9@26_g N_VDD_Mp9@26_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@25 N_OUT9_Mn9@25_d N_OUT8_Mn9@25_g N_VSS_Mn9@25_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@24 N_OUT9_Mn9@24_d N_OUT8_Mn9@24_g N_VSS_Mn9@24_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@25 N_OUT9_Mp9@25_d N_OUT8_Mp9@25_g N_VDD_Mp9@25_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@24 N_OUT9_Mp9@24_d N_OUT8_Mp9@24_g N_VDD_Mp9@24_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@23 N_OUT9_Mn9@23_d N_OUT8_Mn9@23_g N_VSS_Mn9@23_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@22 N_OUT9_Mn9@22_d N_OUT8_Mn9@22_g N_VSS_Mn9@22_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@23 N_OUT9_Mp9@23_d N_OUT8_Mp9@23_g N_VDD_Mp9@23_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@22 N_OUT9_Mp9@22_d N_OUT8_Mp9@22_g N_VDD_Mp9@22_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@21 N_OUT9_Mn9@21_d N_OUT8_Mn9@21_g N_VSS_Mn9@21_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@20 N_OUT9_Mn9@20_d N_OUT8_Mn9@20_g N_VSS_Mn9@20_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@21 N_OUT9_Mp9@21_d N_OUT8_Mp9@21_g N_VDD_Mp9@21_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@20 N_OUT9_Mp9@20_d N_OUT8_Mp9@20_g N_VDD_Mp9@20_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@19 N_OUT9_Mn9@19_d N_OUT8_Mn9@19_g N_VSS_Mn9@19_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@18 N_OUT9_Mn9@18_d N_OUT8_Mn9@18_g N_VSS_Mn9@18_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@19 N_OUT9_Mp9@19_d N_OUT8_Mp9@19_g N_VDD_Mp9@19_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@18 N_OUT9_Mp9@18_d N_OUT8_Mp9@18_g N_VDD_Mp9@18_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@17 N_OUT9_Mn9@17_d N_OUT8_Mn9@17_g N_VSS_Mn9@17_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@16 N_OUT9_Mn9@16_d N_OUT8_Mn9@16_g N_VSS_Mn9@16_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@17 N_OUT9_Mp9@17_d N_OUT8_Mp9@17_g N_VDD_Mp9@17_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@16 N_OUT9_Mp9@16_d N_OUT8_Mp9@16_g N_VDD_Mp9@16_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@15 N_OUT9_Mn9@15_d N_OUT8_Mn9@15_g N_VSS_Mn9@15_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@14 N_OUT9_Mn9@14_d N_OUT8_Mn9@14_g N_VSS_Mn9@14_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@15 N_OUT9_Mp9@15_d N_OUT8_Mp9@15_g N_VDD_Mp9@15_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@14 N_OUT9_Mp9@14_d N_OUT8_Mp9@14_g N_VDD_Mp9@14_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@13 N_OUT9_Mn9@13_d N_OUT8_Mn9@13_g N_VSS_Mn9@13_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@12 N_OUT9_Mn9@12_d N_OUT8_Mn9@12_g N_VSS_Mn9@12_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@13 N_OUT9_Mp9@13_d N_OUT8_Mp9@13_g N_VDD_Mp9@13_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@12 N_OUT9_Mp9@12_d N_OUT8_Mp9@12_g N_VDD_Mp9@12_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@11 N_OUT9_Mn9@11_d N_OUT8_Mn9@11_g N_VSS_Mn9@11_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@10 N_OUT9_Mn9@10_d N_OUT8_Mn9@10_g N_VSS_Mn9@10_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@11 N_OUT9_Mp9@11_d N_OUT8_Mp9@11_g N_VDD_Mp9@11_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@10 N_OUT9_Mp9@10_d N_OUT8_Mp9@10_g N_VDD_Mp9@10_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@9 N_OUT9_Mn9@9_d N_OUT8_Mn9@9_g N_VSS_Mn9@9_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@8 N_OUT9_Mn9@8_d N_OUT8_Mn9@8_g N_VSS_Mn9@8_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@9 N_OUT9_Mp9@9_d N_OUT8_Mp9@9_g N_VDD_Mp9@9_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@8 N_OUT9_Mp9@8_d N_OUT8_Mp9@8_g N_VDD_Mp9@8_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@7 N_OUT9_Mn9@7_d N_OUT8_Mn9@7_g N_VSS_Mn9@7_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@6 N_OUT9_Mn9@6_d N_OUT8_Mn9@6_g N_VSS_Mn9@6_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@7 N_OUT9_Mp9@7_d N_OUT8_Mp9@7_g N_VDD_Mp9@7_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@6 N_OUT9_Mp9@6_d N_OUT8_Mp9@6_g N_VDD_Mp9@6_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@5 N_OUT9_Mn9@5_d N_OUT8_Mn9@5_g N_VSS_Mn9@5_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@4 N_OUT9_Mn9@4_d N_OUT8_Mn9@4_g N_VSS_Mn9@4_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@5 N_OUT9_Mp9@5_d N_OUT8_Mp9@5_g N_VDD_Mp9@5_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@4 N_OUT9_Mp9@4_d N_OUT8_Mp9@4_g N_VDD_Mp9@4_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mn9@3 N_OUT9_Mn9@3_d N_OUT8_Mn9@3_g N_VSS_Mn9@3_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mn9@2 N_OUT9_Mn9@2_d N_OUT8_Mn9@2_g N_VSS_Mn9@2_s N_VSS_Mn7@1159_b N_18
+ L=1.8e-07 W=1.1e-06 AD=2.915e-13 AS=3.1075e-13 PD=5.3e-07 PS=5.65e-07
Mp9@3 N_OUT9_Mp9@3_d N_OUT8_Mp9@3_g N_VDD_Mp9@3_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
Mp9@2 N_OUT9_Mp9@2_d N_OUT8_Mp9@2_g N_VDD_Mp9@2_s N_VDD_Mp9@4995_b P_18
+ L=1.8e-07 W=3.3e-06 AD=8.6625e-13 AS=9.405e-13 PD=5.25e-07 PS=5.7e-07
*
.include "inv_chain2.pex.spi.TOP2.pxi"
*
.ends
*
*
