************************************************************************
* Library Name: Lab1
* Cell Name:    dec
* View Name:    schematic
************************************************************************


.subckt DR vdd vss con1 con2 con3 dec
.param Wn=3u Ln=0.18u 
.param Wp=2u Lp=0.18u 
Mn11   dec con1 node2 node2 n_18 W=Wn L=Ln 
Mn12 node2 con2 node1 node1 n_18 W=Wn L=Ln 
Mn13 node1 con3 Vss Vss n_18 W=Wn L=Ln 
Mp11   dec con1 VDD VDD p_18 W=Wp L=Lp
Mp12   dec con2 VDD VDD p_18 W=Wp L=Lp 
Mp13   dec con3 VDD VDD p_18 W=Wp L=Lp 

*Mn dec node3 Vss Vss n_18 w=1u l=0.18u m=1
*MP dec node3 Vdd Vdd p_18 w=1u l=0.18u m=1
.ends
