************************************************************************
* Library Name: Lab1
* Cell Name:    decorder
* View Name:    schematic
************************************************************************

$$$$$ .subket DR vdd vss con1 con2 con3 dec $$$$$
.include './dec.spi'

.subckt decorder vdd vss con1 con2 con3 dec1 dec2 dec3 dec4 dec5 dec6 dec7 dec8 

.param NW=1u NL=0.18u
.param PW=2u PL=0.18u

*********************************************************
*.subket DR vdd vss con1 con2 con3 dec
X1 vdd vss cont1 cont2 cont3 dec1 DR
X2 vdd vss cont1 cont2 con3 dec2 DR
X3 vdd vss cont1 con2 cont3 dec3 DR
X4 vdd vss cont1 con2 con3 dec4 DR
X5 vdd vss con1 cont2 cont3 dec5 DR
X6 vdd vss con1 cont2 con3 dec6 DR
X7 vdd vss con1 con2 cont3 dec7 DR
X8 vdd vss con1 con2 con3 dec8 DR
***************************************************************
MND1 cont1 con1 Vss Vss n_18 w=NW l=NL m=1
MND2 cont2 con2 Vss Vss n_18 w=NW l=NL m=1
MND3 cont3 con3 Vss Vss n_18 w=NW l=NL m=1
MPD1 cont1 con1 Vdd Vdd p_18 w=PW l=PL m=1
MPD2 cont2 con2 Vdd Vdd p_18 w=PW l=PL m=1
MPD3 cont3 con3 Vdd Vdd p_18 w=PW l=PL m=1
.ends
