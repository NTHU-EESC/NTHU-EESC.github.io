.subckt inverter vin vout vdd vss
Mp Vout Vin Vdd Vdd P_18 w=6.0654um l=0.2um m=1
Mn Vout Vin Vss Vss N_18 w=1.8um l=0.2um m=1
.ends
