*103061129, 103061119
*2017/06/19
*only bw<30M failed
*vdd=1.4 iref=55u

.param P=100 M=90 N=140 O=90 M21_m=5 M22_m=50
+ M31_m=40 M32_m=10 M33_m=100 M34_m=100 MC1=13 MC2=20 MC3=30
+ cm1=10.6p

.subckt  AICopamp iref vdd vinn vinp vocm von vop vss

**BIAS** 
MB4 iref iref vss vss n_18 W=1.2u L=1u m=40
MB3 Vb1 iref vss vss n_18 W=1.2u L=1u m=200
MB1 Vb2 iref vss vss n_18 W=1.2u L=1u m=200
MB2 Vb1 Vb1 vdd vdd p_18 W=1u L=1u m=30
MB0 Vb2 Vb2 vdd vdd p_18 W=1u L=1u m=43

**STAGE I**
MM11 net01 iref vss vss n_18 W=1u L=1u m=200
MM12 net02 vinn net01 vss n_18 W=1u L=0.5u m=P
MM13 net03 vinp net01 vss n_18 W=1u L=0.5u m=P
MM14a net02 Vcmc vdd vdd p_18 W=1u L=1u m=M
MM14b net03 Vcmc vdd vdd p_18 W=1u L=1u m=M
MM15a Von_1 Vb1 net02 net02 p_18 W=1u L=1u m=N
MM15b Vop_1 Vb1 net03 net03 p_18 W=1u L=1u m=N
MM16a Von_1 iref vss vss n_18 W=1.2u L=1u m=O
MM16b Vop_1 iref vss vss n_18 W=1.2u L=1u m=O

**STAGE II**
MM21a Von_2 Vb2 vdd vdd p_18 W=1.2u L=0.8u m=M21_m
MM21b Vop_2 Vb2 vdd vdd p_18 W=1.2u L=0.8u m=M21_m
MM22a Von_2 Von_1 vss vss n_18 W=2.5u L=1u m=M22_m
MM22b Vop_2 Vop_1 vss vss n_18 W=2.5u L=1u m=M22_m

**STAGE III**
MM31a net04 net04 vdd vdd p_18 W=1.2u L=0.8u m=M31_m
MM31b net05 net05 vdd vdd p_18 W=1.2u L=0.8u m=M31_m
MM32a net04 Von_2 vss vss n_18 W=2u L=1u m=M32_m
MM32b net05 Vop_2 vss vss n_18 W=2u L=1u m=M32_m
MM33a Von net04 vdd vdd p_18 W=1.2u L=0.8u m=M33_m
MM33b Vop net05 vdd vdd p_18 W=1.2u L=0.8u m=M33_m
MM34a Von Von_1 vss vss n_18 W=2u L=1u m=M34_m
MM34b Vop Vop_1 vss vss n_18 W=2u L=1u m=M34_m

**COMPENSATION**
MMc1a net06 Vb2 vdd vdd p_18 W=1u L=1u m=MC1
MMc1b net07 Vb2 vdd vdd p_18 W=1u L=1u m=MC1
MMc2a Von_1 vss net06 net06 p_18 W=1.2u L=0.8u m=MC2
MMc2b Vop_1 vss net07 net07 p_18 W=1.2u L=0.8u m=MC2
MMc3a Von_1 iref vss vss n_18 W=2.4u L=1u m=MC3
MMc3b Vop_1 iref vss vss n_18 W=2.4u L=1u m=MC3

CCm1a Von_2 net06 cm1 $[CP]
CCm1b net07 Vop_2 cm1 $[CP]
CCm2a Von net06 3p $[CP]
CCm2b net07 Vop 3p $[CP]

**CMFB**
RR1 Vop net08 15K 
RR2 Von net08 15K 
RR0 net09 Vocm 10K 

MM1 net08 net10 vdd vdd p_18 W=2u L=0.8u m=4
MM2 net10 Vb1 net08 net08 p_18 W=2u L=0.8u m=4
MM3 net10 iref vss vss n_18 W=1.2u L=1u m=8

MM4 net09 net10 vdd vdd p_18 W=2u L=0.8u m=4
MM5 Vcmc Vb1 net09 net09 p_18 W=2u L=0.8u m=4
MM6 Vcmc iref vss vss n_18 W=1.2u L=1u m=8

MM7 net11 Vcmc vdd vdd p_18 W=0.8u L=0.8u m=15
MM8 Vcmc Vb1 net11 net11 p_18 W=1.1u L=0.8u m=15
MM9 Vcmc iref vss vss n_18 W=1.2u L=1u m=20

.ends
